`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Fmxiq5J51BcP5J6at0POFoHSI9nUrlSYILdqUrjuBwVK/YWrc7mQAtfL+F4ZdC2RuEAM0SHYoorg
JSc91pGEkQ==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MLmhMj3JIvJn+WmgTWL9ohm3gRuFd3uZjWtopExvsot7zJ+4eaRBk7mcqQPItokjJA3AmjWAm7fb
lutj1qUXPDR3l25YdRM0suWc3POAil/snJ1rKUdDOviR3B5TxdIgsSl0BvvJuKvz5AiHZ5BITMxU
1St/WyU/YhkZyRTGgCg=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HFRHR5gfIlvfh6z14gwhsBs3aoV7khzFoGsqma/ezG5LdjNRVreY/zBjAQKUjovPWUB7n3N6Ve28
CNMHtEDRUsUeEVFsl3KGrrLduLSekVXhkapt25gP0FIaTSt3dpwyU+oBBgIy7qFmYrwoE/IjC1of
nyTgZzPGGG9evmTqrygBW9UWmXBks/h8YFVLK6TZ3pIe0s6zFWX5uACa54CaWJBIsZ2DjXN3qd/9
aQGZU/xkzzW/V94rtbZF4uYZq8PfEGhTj7hU+l5UdomHmf8FHDizhITDFi7eNtm64XoswVt6u7d3
tXTw+RWK1NvfFDOrA5YNyZB3MJKWIHpweV+WVw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Wm9xIGhssFB3tNW91yRNuqVYWUNmLw67+f/gYna2w0dJqeVkv9iZnLpBC+Vjwnnor9Y4mXxGjOfo
Jobe8xifZT0GsM7I28a/ZglFGFbGUcL9JdkQs5NRCfeOfs7pNUQt6ndMNepuk7F8AIyQzyI2Y9kb
HBbPyhNcxmKcJEATOFqtZ+nMIUsqbMlN3RVm+UIqTA1vxr8ZBr28Wdu+/1f19sUQ6sGSOaLJzCN4
gyLZhnAfLYsgeSplmAaFbY9Nl06JtAcxFJj6DQcptVcIgdLbGFhOaay8S24JYlVig50fIUzUQu+Z
9CgLRge5IdTXAA38idczlOEogDFbgfAk1a5fxA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dua4vGSb2WX7sCjJVXmaQ2+REyd40MD1k/gN84SxP0vnD/ift7ZP5ubkL0Px0XbEpr5wCLYsAHXd
Ol1QzLCwfUbSDUthIcEbu+kvttpyJ59jsYQwqYlOK7Nr2Dl2a7Z3Yys5D2tnKSkg0ai25SFxB5kD
H01v4R278pYhMWkHRPknBHwJZFN23tmRgwafWLdD12rYTT/ch7dWd9oopZVx1lwByNSCjDasZJvv
jVxFNinrlVWJGzQIhmcjV1xFnHEEBuPqCr754lixy/c4q3KO5PUTG5biGIYc3ILdTigavS/ZRsIL
eerN4ZjKO/bU9cxNkXJKKFqpJ/zFO1bmExPqaQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
f8nlZHBRkur4H3IMAFIZTi1PWIxDXT/VH+UucEEaPPmVIAQePmkzBFBuVXb02A3yJzF3ZHpF++6K
6GIL2ATsH6GPTvLd6bmRfSR3hMQLjK/hKhXNGSikMUoIjKZEuk2JBQJTl/RqEr+61x/0tJMHYK42
kEVD3nkIuYuQ83JcrFU=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
F/a2UbIqAwpxXsi0ieidg665Xp3W69cIcPvK4ycZsUlOYfUQjjK6mMrATKZLhnf+zi66iRZ5/CRj
uApIO2OeUe/fUu+FisUAkETCIaiiiSGJJWDHYOphPv4scgmRgCI1AuhX+SWUsMub6CusCYdj5ovL
cDuuf8aurs4FYK0UiEQw4TqJ7nbB7NcmxwmXs9INEtTmtoyU9KsXDH/rRhNQX2MUONRlaFD9OK6K
+b9ynfsGMtA7BMbCq19ZF01rQOGSdDwpJkrlu9+RvM0SGKlesu4vJBMPZjDGN/+E1Sdn4hfhIX66
kmXK98nV4cV+nPlHvSgDTgA1eoGSolnbUzSmqA==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QwouDUuZ/+KXtmCd+GkQkcB9bmv3bXCYGf2+tGl7lqe0qbBqTV3YGqYRyM/D5RMXvryKDOnKN0Eb
MpfbzZ43JE9c2FrZrBI6eJiZwrw6uHhLO3oBeY74IPMmLnhLl3C/FQ0cc+f6lPJ76ofvG9Wp/Mlv
ujd4/6AYp6ZUJmGPT/ojWAWJh5FhyRAikAlxGGmgqAEAkGvMHQkJj6bdpAKliS9KL/2PbTUNKQZ3
dsKrKRK4BfB2Z8D91Ze3TBkXMTFwN8MjapRBSdCXhjjUX3bZBFE8ApF5mkjZjmkMav1+24QdXge5
HlQBl7Z+8uT+ij3A5+q6iRba6PNgEPRGFjTzkw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 566368)
`protect data_block
nJ35GzSPj4/NKoIq7H4mByz3FOcz1VhT5kDGPvDWd1NQDM23heks0cSKEwi4GZSQGkU6PWMyy6CM
TG07RSUiM5XmeA2n+UqZoLT+HskmaPQ9lHl2H0oLoMKGlbnOPacX+4Ia1lM59aMyAwDN2J8EPKoS
8yPrlshGJy6fzx/ffstev93PE7mt2D67MBmehWWAiFFSViUfV/V2ldp4ZWdaJwpvzoAXDbvP7Eu6
3Oul+NNH4uQYoITkKH63/5WvMOpDXWoeC7yOT7FCd4PMI7hHX/u+2GjM1af/ohzcvhwoRrXeLltR
fUDd1IWvIfLzKTBID2gogc1r8G27t5Cqkby5gqyrNB3s29nk41DtgQZWS5l5/thmYSPXE81wyEgz
YNFBt2+bsemxKYCM13EfkBVztKaQGVwj5bvd/4GJKfPY5WR7T0/+BwjngnSffgQZlnoMW+bewYjp
YItbU5qBSzfDT/5K1SqdHkT7dAzDQ5s72GbS5IXYZdFJaHSMDijiL/VHCuiassDv5KFbjDcL2i3a
DmIxOvZbcaN0KJ4w0KiNjbAngu4Ahr8ALAH/feh4e/jGwetf8J5dMKYS98/HHqLDiSl/RRsFibzy
AppgXVoU62GHwK3UXs+y75sg6DWspyHgGRJxl4MG36vlZudT38LZTTVFcRLG/UTKOpLvbxCKaUva
PQKhbdH0exdfBbuazhYy88nMTPG4pQzCW1x6tiWeBQNCjyJVmScwtQhYNoYydu3XK76Rd+XvgVpu
Ucw9xTZbEoaBDN4HIk3HIzTgANtwT7aWWgYFczk8FBdNhNDoNHUoHtDoHiOdp7HzfwoIZK9eP1tF
853tVtgRx6ruA7Se4FJXRy7HeQT/KkJnp33ydknERlzpA2jgGQbOSZ0QoOQINNZCaq6jzwiyY5O8
LPtbrPuAHXqTw8eWbnidtCz7Qx+dxcwbgJY0fTw5tvLlq6MNHNy8BokAqHLEfL735Dhr8KopOnIT
RLI0x9kXoDaCYPu/JPWHYNYfGGn+8I+RZmRdFJflNlQ//cehhHOn/uR2uEgCYrt70NAHD5hpj5lT
9CDhSarEo7tyIyNA5yES6wM3+bK39tOvORJFCY0v7hNy0tjwMhKKazlHqQxUwPio0QUKgBB5desK
pLXep2fTBhmu/ZFq+Jf92PWFt3Jtc6VSaTlVM670c0+g0h9lfDxjTCTESOGB56qc/TDrEM4NMf6Q
YUANm/nQzEhxIzFutTLRDTHTPoQErnQ17GbfvINxQ0RGsXp/zy3ugZqYABUICYm3X2u+1909caWW
9SDTdy2vN++xypH7EeJp2kSfk8uepGjiLr3/7fsO3YtP1gxZFk7d1sJeHcmoS7lNnoaQwiuMC2M2
uQlRLl0nmg7wNem3vn6eCPx0dkSa0cVRmkHhfqIkJjKCjCEMiDH0Gf1sRycAQHyYFa8Ryu3etcWQ
HRH7sgN8QVwnM+ff+UTaN1rVINGDmQnhXBxBGuuS0SpqPS/MCmxU2ZcZ/oIMR2nGyH/UTrYNG4Am
J8EgntR9ELwtIRYAV284q3FLkJQWc5nkZDrnhNukbj0p5uvvYhnu/Z+yo7lwy6s0ohaAhgIsrdy6
fFL7Glgz9h6JVh6APSxgJljKKgMPgeYpxdTITfgXwy6n5adKmRIerXcsfELhbkV3h3AmsetvvKLu
P+UbnLWlXNEKUAP9OgI9MWpiHB6bFTg8EYuUAce51gSfbTDGJhbiB3tNm2jpsZ/t5Xpd6abWK9GA
b2E3bq5/ctKmdxgAZcKmfPKttUERas16xCxmDLGfuYqRrUWz2bZXY9a6ENLEQmkd02Pqxdxutlux
S4cb9aZHrYIguK14E+jzblgYdb5zUrrmcDDhTS3A4YMMSeC2fC7qJrMgLl6URybhunqCqkA8CA4R
KOc7W5nMTrRXSopK6ml/cDcpWXgblu/iNtKNUTcCZu/Zhg/6DysYI++vvtiuTsOG0S47DbxYJkZS
4Pnm/aoM04dj3aoVy6JPzr/Tcj/nmiHlraLmPx7pJFMGWYAW9Tm4HtBeythPOIMzdRUitd2Y797+
6FZctP4veKIkqWjHnE6BPUvMZt/+XGtYw4TmOxw1H3gLgZFeyzg7N2okQi9iRgs6dxaS99AXFpmZ
A790a5R4JT/KhcKNMmS7NTQP6TY2nSamsBu3wQ7ihmbmAxsRPNQuUlOLle2+6Bwsfwd1g9pLlB+5
gEspBygsBj0FTDGJrPEaqnwUppSdIrNFdmFc7C3VSwiePMhYfjFjczx8nZApdtdEfXchuIXYcwMM
J0irTXmKRy95rV0IDT/G98hLsnn5nKcRyYjGqM5B+97IqP4yvxE7kAL4xsCUupBcRfs8vxLALPX0
74m6zyQusum+ExkqxhHkedtk0npAq20VW4vktymgfQ5lNjcQzBmT6IKurv2L5q4BbJ0crxc8bXoc
DFjC0i1BxjR0GOVRvh2RdPp1ojeQIVmW/Brud3Fsqro2qGsbpHN7CMdgBk5AUDmWzO7fszFWJ0nu
6WRXxobpW1+tIwMlAzv5QcQ6Av2Yay1dr5XOJJL5unuNcOiQbATVbVO9QYZhQpeB6E1y6tlegz1M
hI7hcp/KaSax53q/0Ies4/UkJTXeArAQpuCgErfrbA3y/MzbE/OlaOt3djemU6ctWl35iZLEiBZR
c5l3PcWcwmzlJ5eIe4/QzSjC6xHdOyQVaH5D4iJin3DnEeRGCuq9Yr7/QLfeyYVYXOcBg4uzNaDu
Cao4gAIjm4VWY5XGqASa2Y15IcI05d336Ryai3Yjv5Az+847nzuwZnxsjoe5K4IbrgtAJhE0/Q3j
QKd8fXeX/4MpGBIDpp2ENya6zluA2MO2I4I2ADGWtiKpJzXk1xbhy4A+QenJxKlioGkId7WQ0LtJ
HDDWgo9lRwJ4u/BxpNahhUKrlM5mYUaJxvY/hZEiJaaoKvgtc8jruQ6yRBbKuFEtegvs7I+64O/D
8TnUcSwHYoifwkEPUFpky8V2+2bGiwCeOZ6RMxivoajDJgs8ZJCo7l8v1agXfO9qK8Pt4H3hPSk5
M/2CuEmZqkUtko3Dj46K07aNBvfjzWZ7bILdzS6TkK9zq0WngWYSnQaH/uNO9kyEgVCPyYmAW6Zh
fuhakB2t/gUEcUlI+aGMF/g9ZcB52ZC/VuiOdI9JWxwiONu2WLBVDNHC58JKpBcwV8xc5O3E5IiD
3mlQjAa6mbBXw4YoljIAhnQDQze4qQM77i/ijP38RlkzX+gjLhMhQbAYzoWCr6DkfY2x03YvRYhg
FcKargHPMfXviZbfNyG2PudNfGiW/EbQpCnpOKvx2F15uROBANYcVyaiKfMdIsj63cisFkPVM9n8
tl7i+3uL4dOgepk2NbFrQDbDtpCQKYcuE4YbL0MaN7qGFfRmu02Edqf07xddTjI8nBufSsRqpEoZ
Co86AEsO9iRLO0ymko507JygkIxW0UXJPpF8MBHblQCZMMeA15I4bsFWCmpWes7isdo3OylIBEy4
NeielzopSB7o2MNogVPrEkdSZC8J9150qM8SlBhh6Fvm9H5SW4fmQj/3xC0O5AogrGDF5Sey8aE+
ITm9ly75a4F9EenW0d/JQX7dy1HoGbUeczq7VwqWAVNHXm/cwbr+nqpooVYjzeTY85aNoMaoEb01
ZYfAMcc/AC/7nEaIc2Km+lj6Wo+BsHbkfrwhIadZ11fwBjsIf1xf/2jeVXJ1OgvQwlHte5IkmAHp
BWKRKcuDNBNPxR7DBEg82nuWpgJCRZvrJ2ObpTWfhy7zJOk79+CqWB/B92CriQGOsemFi/GhyXwv
3pyzblL1cr2Cv04osZa6m+zmYptQNt0i/ET8+SFLEu/d1Vg5oqHriO7Kn4vCLIbnbAcZTV833BXU
0Xrh/9q36RwYK9UIyUmhaYUa/ChCbUfzvB49TGE9nnDYBoJ1r6dNfk2KMgnYHnlZRExVAEe4dlnG
F92/v+/PtuedI4i/oxJ3N8wYEjAT5hcBIU6y+DNXNEvCWV+nzT7r5YPlWZ6TmrovE6hGjSCmi9rR
N/DYFX5XQ/MJEZei2faX5OUKffOFuw6E4MP+WWTURgumNAQUIMwQ985hjXaCNEwGahqZApy07jMM
ARkEwANxyh084vg5THcAkvx3oc4HZQlyAMOMHg4KYLvY8v9AyMj95bRgnhQXX8Sl9cWf2d8FB+m6
1oPOL1RsIxSDsEy9uRaEtMZE0jx4U8SP2EOPPcZQXZo8osGFABWW6b0F3e2pe+ay3cvdUglChL1l
1HGyFyl5BVbnzN4zifXKNuCq87IoltQ3jeRRB3X8t+JisdYUMTEC5B/9+gUqIHzLrnzQl6px5GuG
wX/hJXLyp1iikcYJOh8D47UaWd5+q7Df7mCoNzce+H7valrapy4dXZ0e1ex4RaEYgu2eMLI7N0e/
wVuJgGGVX3Z4S4yXRUryfFzwtNlLMdlbAPHKktpY8CAG86tA0yus5Egelop+iLpvC8zTHQFjMyN1
kpxjSI1SCaj0TOx22oSp/CGSfdYDVd5B0qdJQxh2NnwuWeiM1dJjmPtO9qVq5f5ret2AoZ/mZAOH
Jz0PvsdINwU6C2RqjEScYw+yeRM2XrqIYlLvwRuGVBdnqLxI0d4i4yp/Hazzy+GUsnE/W/oQWBmn
QcSMjdGgVHr7Oyqza2xAzyJLAJNyb4fVBupJELSlVR6xKhWeFWOj5nRxltfWIZBwokhDg6qkU+Qn
vGBrTU3OFYLVZ1ogcTEPdqCtnhg82P0P6Ob6SLriMgJpsVw0j+C43OSrTdOD/1pHpkzcwFZVhun7
/pl/Aup/M6RE8FQm4FWmFL60fgd8gZdZ8tzcRaz2HlxYToGtlNKKWj0wyOWgWxDk3FaOxAc4EYPf
lqqGpK2nCkijc+DDusigpncsnVQeLLsiF5eRY0fYr6yX+OSThJkGGWaAwcyejQfqsw6frduzI9+U
P5y2cAiqs8L4ohW88K8rzweOejeM6w0eCO6k27jrlFpMewO1MHklfK7rf4sfHdABpaSNpqsGTayM
OXVJRo7H+RVKT1gCZ8o74il9vadT3smHpjtkGPPT6bk68eZY9zKqDp3PzDOeUPAv3kqn1csKZTTJ
V2JD23MTwaQgJi4vICpYDun/WEKL6/VvnAUkvVFflkpLBJeS4d00l+23Zkhw/2Nmi7rxfi2rpPU9
F9hlPStbfwJUC3zr/L3mV9FyfDlvcuxt6giIv6PiVmTDxMky+Vlt6lYdn4gxf2jeDhVbecP3DiYv
MjEVfhSS8TSpUVjHQbLxEWH7bK9Eca/0SelBW1XYskEQYN5oHJnhMuE0Vc9oXWplC+0SO0G478hO
gPn/l0gl/FP2l8c0cCQUhSqlTeOPCgXIfr6Mq1YpawIm+8ztmhYp72cbzAAtOUTDypZAYi9lHA1L
za/kjaHGQL3TmBf4EDO7/+MzkwQNBh8Li6CNp3NqXcs/hlN8vAjFycQ1rqqi5WZ6S1Rie2YZ6PSj
hjMuBfTeQsfClI5qvORpKH1+oE+1UxGVEqbIQsIXO6qUQh7B3sp0RVr7+NEsbxfwIuIKwRDeXlty
hXFQlQYiz9rQMIB6M9u1kUmyXyJ6EaNxGOZ50n+PzWlfSgBG4X4V0Vg4GmZa9Iu6aTVxAIsW3a31
SuBN9ILjfjYmDvqe6UK85wNRUZKKmwLWQ0ccEeDSCh0Es8rUJP0DgJjlleDEU1DTNpWUM6fZON8z
PFnAFTyy2OJTu/UDHPkTe4l7f4uDiy373y4hpJXkzypJzbpezG8oKwJ8jq+BzDRRhQjRS89A60HT
37QhXC5GwTVm5/x0Mu+QTCDxe+Whj/N89By6cT+HqsHeqaeyPD+nfgCtyKK0V5wEcLB05zTZuNxw
mGdBaUCxUTgNGDotXNN8x7OUOzmZMm8yTIvGlcDUvRZuQc+e0syfmdaWYDOHjXk8WgcriTHR39Gt
zMtfVgfj0Kt8l3cWPpBGaKSJ3vv6bR+igsFP18rTThgtBLXLswRQm5i1OkirEtT2fpl/38BpWbYp
MBLhpTXDt+fhE+Jk6Q9ezW7DELtwFV4zKmaRhUZqPeC7eA0ZPz2RxJkVJ6Wxlny/OayW+BfdAGHx
+bxwEoAfkTc2zdQV4LD7WNIDqcdvrX4HC3U1mWWLqWUxKo7s/02zY8Gc3/i4IqKBtxKlbsKhsFT0
xEaZRAYr+s8JHJT86Ch7INEXHgWYqV5r+EkZ0ZJv1NIRXfryq2qS8S1xh3OvoeLywei+ksRt/pss
Lb0sYkR28rB5T7njmCp24Dz+XCmyjBinHc6+wUGpAGxWNeemvaiw8wn1/EPFAmezIaHm6+0DG/Nc
tOeh1a0YqqRLWqq8huE779P+iLma7aB/8vfOn5hdJT7HutZLcYE+t2F6bffUpacD93VFz6W8OLYl
snUO40Lg0JZpfcbqjyuSy0PiwibJkH9bRnL+LOUvkS/vAmd3swDOdVacljJ+STFtxkkabqaaD9L2
4dvRbhjs5R5VcKjw6vzB6CmDX1HSo56V2eJ7bKR3zGOy7ci/6y/it6M6Os3T0dUnD+6kFWKj+1KS
1w4ye3kNXjQ0yu3ATFNvZweOIuNPYmbCTqRS787Tedp8VOYlZ+GYLVEWlMxk8XMhb2asyp5BV9cZ
7WisV9s67qLiVJvN3JQeKl0SKdkBEv48oTxhzN8gvHPlHGtVXwVrlbi3HXYU46qw3QBBCBCtvzvY
NQCvziwamjkU8IScfEylQDpYLc0XOeEtY6/sBHxW+B+3DhIKUKSoeeORtxpf7CQMqYbl+K2BhDIX
G3Neyvn0Hr6vhAcehTlTYPfOvJzg4QfZm+hEr7eUa13eUFOFxBNauOBzN8tzChW89AraBQburdN5
X0VN/755v1IxyCqsrVj4LbNRWOoJ93Jh5nhoDGgbuOeoXfZVFNXT76JObLOGNnhaebMKXWjlzqQR
A/5SGO6NJOocBCmwZR9bqYAJOAMrjCXD5a1+j3iIaabemEsBmweVlW2X0FVnWg3GeCo+YqFW4eJH
+ehC91ay+/Hu8ZAlVZi3WtkjR8ZK3zdyKN4dSSk0pYa/JIz6x3Y+A0h8fWmTybdkgk6k9qyhs5MO
HdTiK4uTUww8INIuqriDSu5v/mxIfXIpxdSgsfSY6AQg7fojtuZkf+PScEL9NvdTgrMEnTJuuqD2
bLpJJ/sUh3DIr0WTQ/WzzzT9bu9dhBS4nHex/bP2ZnuR2J67+p4UuIYKQHwj7TqcRfsBQSs1lR4g
uO1a+4wZdc84+PschoXmLcvNSZf2VolomjtgtgVHkbNuTtW9RgCm0u+H+480ET4MTYHN//f/TJQF
Yja1rR2HWFe0LjwSg5AILfXIvdNCPyM53ZpUgWNjDBNKi/rfvjZ8xYIOV6KhTOcSmvEwiEnE2ymO
RqkTV+B5YwsUr/MhTBzGW53b0Q/fykkeFIovgmulkEuANnBwlF0NldJw8+s+Vl7KdWCU1EAruUCq
XicBXGJSpGj1ktW+HY3raDj9pwafgnSYMcQ37uLBT89jd9MhsI3bgPsvy0yPtbG6mNxrNGJKO6o8
wPmyQsFOmPJ1CJAgshVyuQfSGloDlKYnv5buQEOYb42qJpzlDsRj1JyBRa/WvfcC60VwiItz2a+K
TY8ycPmBjHj5wXcCNeteti5wvICUY2sdZ/QPTmvzt5bgLeTcoFrsB9PvijIyaZq1rK7KZ4vlauOq
mh0k6ZzmZpQa7NeRYMaL7AUyZNg4aMw3Ezwn7b8Mh5BJF57wtbW+3t3uMU85SAN3SBfTdPukJjYK
7znS3Vp8vsJ/JVJKqMbEJIAnx2iMoT3w0rN5PGPwhp86pOynSDGoh+o/6dyJu/Sg/THKNoiDaQcn
VFgNkqNCgqWd8+3TlQxDqeYDMy3Kllp3thKXSomrFAW2h11hUThP4DnWqLlGawF9Q7XyL6OfVrWb
UEn1etZxVVw4J36Qr+3nfg2oXFwTlumYjwq6nceIBf3UAiTpuqZ4BThq419WLwyK9OLbWIq82ScN
Jvi0LLQ4FUYxFWvGiuf/UYQEQBRADpwRto+EmOL1cT6x3y8PUtnktkuXh+vRKBkoUIE1D82uZIfj
KXuYn+GGm1PqUwCyd5iy6sLI/icf/wnr8XZTIVZYdr/t06wS1FgQghSrPOjxX3m8FkPRFCBq6mET
Tz6vXrZI3QT3WLUPxt+nCh1FWdJ0Hf8nFWkF2XC9wRR/swerjlITeM8Za692UkXDyP7Dfak0KBTv
lrqab2aDO2ZQr7f5hYqWm36dRxPrLGoOxL9QRR2UNw2G3Ow37gnZGHk09vnPqe79qHHOWFCJ+vdL
HN8aHaeco0XPqzWGYC5EEgnpVRIIRADCWctBYWT69YysE2vXUKhpiwOWVB5g4z9GADLVhYl/EGxW
NH8gIC66yl0cEwVAAG0v+NLQCtP+VNg9n/98rDWfZ3syax65hxgCpbXdcxN82ZsRT9FBCaX+mS70
zl2Jw8PLxnKsunixFVW+anUQ9eftap+3/DFrsAK8kCzrT925VPHcIfIKDpyM6qFgzJCrH34jILC7
WjWxe2GCb/WYqvYmaPUqa1MSacsE5ndLMnuqYAUzgaaSbK6GalVX3PUZGNxne6o7HpjIc+JKQyew
Lu6eRtBNOPKHZDxDUr4dHi64E897W0NqQU1J7cDoD6QOUeaIq+5vQ3qHk2sNOUG5AwlNpmodcOgk
UUWCYqU77zB4GXpt1m0k9TQmEPnSjqOUDWQAgf7HdBiXjLiG2y028qWRzxoPX8gNDakd5XikH2Dq
84P+9855qsH7S/2BEsSbcK5m2ZDlE2YeoLGfp1JWF5WuFm+YzkJSRZJz1n0XotLlaZbKd/8rWrqo
CUuVqGfnat9JzxrH8wCGN7aItNnGnGtmv5Go7sXTrVlHKVetiuPYNXRv8aHRWgFlnagLI0vmcx+z
xSzClqOOBXPnRNqu5yUW7LXcPRRiSGk1l6DPNv8o5kqPfs/ZXTHdOutB42I+fOpa2Xj8N9hO3zJt
nvCvhl0Rli2RwTs0gS4v7e67GIDfstcv/Y8Fi387Ge+COfjHrv3CsBxe/OhCbGLACCQ+wSgw3lLt
E2gRXBKJxZRZMH3c4Liu3Zg8zps9p3M2N7k6EBknvYsj5wFBUkBzNLwxNYttE4BHGkhoqaO70/De
0ZhANH1x68lYpweGXUm86YlyMsII7cZcCBJWQwOFR6QzuFdtSZIrJPZFZJlcC0MrsI9yBpwTLFyw
/CfKCbQ5MLkOPBmrXIFA/apUwx7lZMq45StB44jeOI9xNVHWsGhJycT49HglEDKQBQJQIRM4RH7x
AKJ88TBl9Ce8bmsvjeHY2t+8Qjiv488szzCQboG4wTGPrGssMz1RiDtQRP1cp/l67EwX96EZ07gE
BujpPabpfjCNYEiJML1FUcrZpLDYADZR8/3IlrTaZ96tMIC/iL6A9mqfJfDcbQQJrXAVNhQgC6eA
AQN4TrIVzRL0KmevCcZbRv8cX1uyi3Cy529IC/RLpbDJ6r3fUxLRfgDrSmYG/r2/3ScxJfSmMIPt
BD4X9yC3NvFAOgndJwZth9wPd2OPJqBhTdvMGPlYXROj6EMM+V093gzu5J2ZLtvq8qirKyj+dlz4
h1BG68nSg/THVAW1gDTRtzd9i8OxVCBTnmH9B9TE10WfJY3rx/+d8bYJNojfwFj7bEBDmPh1h89P
7EGfIoarQkkMlVQGcljhywAUAm+LSEBH/n3R/zmjHXgYJCUeAvjh76EbsT4p+DjvO198S7jdix8Z
bqYc2+FOu3t9lDfZ32xDN4PMs0rfZ4tAl39Bnx2Z2fdQ2MjfjdgJJ85cr5Cbh5yiZFcvr2wUhu1/
g+7RfQkEi3sKf3hM6b7Ti4vW13IepFsOVQ3cH20CQOhWTBqqjI6bwR1SqO82ETEyXYKEtSKFjAm3
r707ZS10dpoqmlULSfAf7hX0dKBCKgjqPTMPuEcylhfKX2hrzmWZvVq0G4mrBLuqFWDnB+58ZIFy
tF4b3/WR7InHd1GmypEGFFe/WymzM9YlYteODJjjFkRaTAwds4UFIMxJyn25Qh3HpFEY+t9/LBa9
BQYgySY11swo/NYDUdL9GbAVTOA1xXTMiEoCq8FJD9v4yqqbbmkEkllG+iIph/9iRVfdfAcIeyKh
14QsmmamhGKFlWUny+Hjlj7wNjSF48VjDRY0P0yIGUpFZkn20xeVKa6u5DbZnGxULucta/U4J8Te
Suwc2IZ8KPw1mzVnZnl/3dGZ3iuyH6UeN6rUNMQntITpfhg3DNWlvnGLAcVsB0gRLx1zwGdiS0YF
344mW83WwIXE6KKari+BjNWkuJUx7t+nVDeDkk8ZvXZlM/I/QgRPOggOImW5xNtSJACF3O25uLz+
j8ZfnW5Vb7BWwMHk0iQPjjyMob86alWfYwzQdUsiPThGkQwB8epcRGQTvE6def9vmkmU2KjLXGI+
Q62dnlhO072ULETfG1i/J8qPbCfkRN49ZbFNQlmGWH5yxXMJI/eVHjcsCBwyP8O1JfQt3BuwMyNj
rOQwtcBi+KpGZ2Jk8Is6AfjhWWxR56N9RohB1Br6+XColar2FfzfXAlEM75S23YoZ04j5Q4Ux5XY
zGyWXPBGu9LAgSf77v1KdevXZEVK4+XeKlfazvf6L/KQJfOw1j/YuwNFXVB/nHKBPA4CCVAVOMr5
Zddt4RsoG9QKnhiiMD8SkaMGOqaKsUsIwWsYhUvsvqzt9vfmV5XsONqoBAwWc7WuL4spTM2ke7AJ
yz/3U9RniOcLpZ4rYF9mBQjhl7Q8cM8HVvua75btkiKq0hA9zd0XjTQyNKtDZo8KF2b2kcgaAWnw
9mVb8J0moXpbd9Vbp0RBtSvFFylYMvR4d6WbSsQ57MVJ4gMz5COgcxCHiFUpxtVYT4nJhDHZbNWF
ohySKTbGqhAONt1QBlea7fnOvcXpOVUA5hu+q5UEnblEh9d18HK2r/jy/SkWZmWvjSo4oFPbMZAr
7SDKoQ53Ncd5rYE7dXh3OXbroclhcpG8l777q8w7NITDVoBSKVtVF0y0vtNAUlQhkjPMcVf1Jw8G
/S5eM+g8fXLfmEAvjhSFVhX/DwEBVqV5lf4/eHbsZBDBr3eQ49kY9/yyNSz47vP2zMxyGkmgkbad
X3+/nYpOuH9sFRz7p70ncOnO0zhSLOFnxJHJoOE492urTjt1kOdaeAhbCmXDT922FckheRRVG5qZ
qEda/A+Ka+kDA7pimAlNi5ZLdothdr0b2pxzRaAbKsu7lv3wpNpTyrfwbD3AhxMZHFWp5u1/FE7R
ujGcONv9EROa/peT3DD4KgQDDXsqVxH6/yTwHwv6S3YYnMvrHXJaBjdFhTKE2cm/QHEkwVXpTgtq
GHyhMBF06qCB9y6XTua7D8zYHXZRnsuNKrg82b9wyvDZsNSx0CvC7KbzZ33HhorQhsPhHxA+//PO
wpR2eEEBWOb32tuDwCZJS7gZkr1rF5yj5ypA44vl8wt546/kDPkjtauXuDD46bSX15FrWr/xGsxf
v+FvniS4ZDomKd3jGTgzyFrRETrRr6iHdm1i3CTw6d13CPF/UGxp4WUT0H6ca/kdFcq+HryhFPjQ
ojmmo5IzgeJjPV1skVcVKtGrlBBtBVW0bxzlE4VtwZrVWjAMtYLrl1Q7/ZJUJl3cLJCUrLWOJkRC
7Qwo8CRe1VgpKGFZt8CeBAp5CCeUZU+HII2gX3cH8QL7qKI2rSWW1dpOTe0s/e4dXR650GMRQ6Hg
hi+awcfM/dZUy9vUMaM0gH/Bgg033GiWOmeiPJlhqLM0o2v1E4Od/w53D3qdnGrPiZp1nGnftSJ9
rex4FAHv90F+ZiZ5QCXuf1uQjJ6kNd9GgmRPxgw8RCBIKpgSAcm7uG5lKoT28+1oQntwNLZYax75
1UCjIlCMtT7M0r8TQYPkUcFC60mwisqm89jXw4JBPxHMpE7tte022oRLiQggv95ZU3yDKzPpRclm
fGBPGIW2C3WvsBox2yf9Cds6aosHMZWLdFr0U2ImBf9/SbnsK8xEVMy6ARJoG0ZDaBt9Yg/PywJq
yhXe4HwPDd3j+CDUYVwkXTScyVNm4WjWpFSCYqj+oKeoj7KvhMKRXDV/d+pu9oBoDUlA/GNYhVzX
xAfMrkRNnTOlblrU5JiThgcq2qa9vGIWQPNYXPiOhTwhMOKFHTAI/klyahp5D0XAvHbl/Hx27Nxq
giFsmzacFJP/nlUgG4JqYg544DdmTN/p2wSpzNcR8cn6xiBDgzfDhlSLh//34+WcJXttq6sqzdhI
gMUsjf7MTlF1VQ2IAAUv3CQhDFlVChjf8p6txvpvCmf7gvYGNmfHhUfOqb2QFmujv8x6mfkln4iU
/5B7GaS2U/L4fIMtCNPOWkJ/H1XHI6o6ge0+xA+YE3pNfTrIgpKfw8UgdkVDz7oluaeduBKoyv8e
Re5Pgvwe1E2I0MbSB5jBCBhVa/gGLANGMavhPclMR1k5SpfzaRGbtMTyGIIupsvW3IgMRJ+Qxy7w
mYh86e0KUqMJETMP2LOsRlwWPfmEPAlU8cVuTzmIGCEPuQeWxsi0esh6yz8wTfExQleAesnvmltr
TJfIDzdSlMbe1Ydvo0PBVAqb6DlO28C87kXMcCKPYqCQAjUu//RoiwXyThcZm3llhGmZgUvmxGe3
i5xe4mYdAdAoZIVLvJ+NfGs6b4Z9g5Gq3DVsvzgyzWDzYQjTaDg/smzRk9YE12hOeTd/CE3RawY/
KB2hzzQyOlXKX6CDEHzM07+l19v+SQgpFx8IW9hKeUNaBNZCR0kE1inGC5Ous0k48+2p8h6bIqE+
PhXbiQZZdQLOXqXJaoBAbrduw6/7hwuSt6GFTzB7K3swX5wFcFGl3IQ68F+x0ueawFWCZVxAtlOI
lLkquoVSweVeCGN7v/UX6xFUFCSEomyIq6a6xNDLefaZdSMJ/K7wiDIgJ0ilr/m7jIe3C1p9Wf+Z
DqIKBm++VD+9RSA45O732jTwOnIZzmvpFWL3VTe1TIKigFL2wC/OaOl1WDDw+dPcreu6kQ3lCPrC
ly2mArHBYvHW3SUQXTvTAYV9Bv3m9xNbQI6bKO8GthIvBLZl5z5ZX3LowtWa0Oq81e9larIpIdLu
yPLY6JHn6dOTfq7rp9KXgOFC5uSMsoVdnTWmeteWn1c8NJyIo/AdpsiXnoYmHmzb9UXTo7El5jyg
qTeQCfCSnvJN3F8E1vxFYKFiFvnTzQjyA0SOgx+lCeZGoFv+rHGJmAuVZ5jf2Q/tfPVWsDEMMw+A
i+P5daPz1T6pFixjebfsYdjInjivU1QRrAwO4ge7h278TPaMYI91Kd2W5xubZcPnDLvyA8zSYMQ3
zzJTSLVS/uPwIgp7iSEdXCdAiOeF6OeGjd1Z3imO0R4J/Hc3yUkZ1XPlzr9xeTRlFFoVCcD5AN5X
JOdKkhDeefN7eCuAWDt0LOX8cEhBjNeQMUBFVCfUEH7L444BcF7Qh1xoIz5bhYKr2uUkpjWNtjpC
om+7pWTpBTzPjZ4NLgyAlWwJ4cJtG2YhnhgB9bzDu8mCuMxwxeX6lopvnObG0iKFU571dbXUlm8S
byDKJfTMYhjxz4skS7+5W3Cp+mCkxfWt6lO7gZa/G359pOqDt9mtPDIZ6xXCTZ8NvkKsAZcioS1M
DUt//7lUhohYw+LGToUePTQYUtYRSlrYAun5Dil/6t/8dk2XyCUibee2v4ZKtvGhqKtTxbLNMxX5
eT6Tw/nMLfUoAohKxeC2lAEOGmpqvI7B9suA7X9w90jJYHu8tt1+r3Lt8lUdwcgn01IxFq3G46yQ
oGuKCyFDglWtgFuBfGHqFZy9OpK7EYHihM1rhEuLTC/J2FhGwJPd/6xr6L8BtXowF6csRPjcivlk
dow1XtOr6RZbkkvKnRfyh3KOXFTnSQ7IirmxGEbzq00ogkWGzG9c2ps92gTUXbSadG0Wil6PgJvV
G3tEagPczLGPYlvRqAHKcUQ8xlrI6KcP5edsDpqQbFokfJ6IDPiHNDsSNtGiD80/x991a/C5YJpH
IuJ6Xtuscz+pg0D061H8g1U6+MerRRaBz919wn8qbKIs060tQ6Yb3GNp0Ge81eOfqtv8r2axlFVF
+83JStsiCXDxCdZymY2w7nL4uu7IpApV8HEHFWbTKsDSt9UlMsco4wqQr2IxxXW6KMjpn31qzXYM
RWfx+kbawSqGxLsb3jkNLnhg76WF+wpkcM8iZObqFbZvt1lBiVDAeGnFgxutHhvtH64TVuRnG34O
smRF8qkusMIRJcAdARkdEtH+oNYtld/mQWRhYoLILyaZmRBhcJWVjCZaQouJTvxIYQ5nk3poH4cM
bJHZ1/lotgGXWpZs9nXk7xbIU4Xx7vsaWke+f1fzy5ff4C+rlClGdZ49iunMyg+515tdQzxhhaBi
ERUs/mjTuPl5pkO6cBVk1+Ph/P6xMaTvyEmEcpJZ+6ZauLy3xqkW1P5BdQoFDyOXDmxpXKVYFcx+
Ui6PEfvGJ6Yz2I4jyDUbk2AJpmoIP8yBX0MY6zptD1u3GrQFekLei6fp2epm31OeYJEfZj1t967Y
72yJa1GVu4Iyst7mzBoUtIVHoAKAPuXYiqHwyPn04yc0B1np9qBW0lfAVeru0bTPhLIUETmo87Xj
eT27et5haJcbniSAz2W4uLJTRutupHEIN67KRR9oW7lZtTGHsjSPA6V/fEf3OsbGuphp7cM+lpLl
DOQdMou10xK5R7wl2/2W/ZJw7n2atz4EE7Tuy6vnaF+rok6btyK5S4ZCYZOWRnVjq+QifvR4Fsgd
uZbKKt7d/g2tra8QVlDo1pzuxDcXnuQRcE9ts0YxlG11ItK+oMsnLcDIF8k/nzNGBGd0wx/S7eAA
E8RO/wSTkOtPZrN9apbtt0y6bTSpjOr5XS2wflCkjViDOsZBRaseOXX2zbjcRbpjD0p3ioZ1JLds
Apjn8eX4D9pMJOsL6vyORInkovPAB4U6p1fWJFV+9Z4g8y3Vtvq6l17n7G7k2g7aRJJXxrrcaoOA
rcB/ORaf5yxCL5fYZC+75fwy1TWmEpjUtW+tID/I8AmzxnmpBS7paCAf06zAcXQMYZGk9QUKBfb4
jCYWvqx8C5dDc6+VH6Cs5feBlCZkk3ccZVvYPvageo8GHYgtRrwzAEH012Fj7C+z0fHQI3u3OmD8
jqjbUKUXR/HoC0GrIpv2civhU70EbTsDT3bqXhzdHkvgGXUwrPQs9ZQkXIY79+q0Ep590OeF0u+7
bUYghSWk9hkOQgNt0oBQoEGflEfUiQB2qXZMe8m89V51cSCUyvPFTaVCagf3DhEyyVw7mGtxBR+m
UlnKsWlR20438ZilKkzO4k21ldrlcbe+jS1E1RhKW3DAYhKzds0iF6YRrilQqAXlEMa9VBW66UhL
8gw8bHk9t1YdyWa476DBO+hfSvbJiPS0WPD47at+ao6f8H7hbrR1Gba4Gq7772+zhdSyny9N/6vt
o2nJ/vSPccoC/c0kz+Bosb3PYHjaFbvgwqywV1YdRYaca7wMjXZL4jLza3w8hL0lKupCLNpd4W8W
1lZwl7JNycppGCjzWOyS+FaMY2iiA7j/FN+hjuP9r4F0sEDbzdgPD0B0qlWvlTyLkhXnURC1KJ9b
qxMUjHzjjP6n3BrOACYP3uGmhv4+3Y3Pdr5rX1bPOoOVIwfp7UqmEjEvGme/sKmmTIamrNkmLq8f
NA6Ux7oJNpF0uoZmq1iPz384WAA/DolOZjRG/DMqh0ypgPY9530KbQuqSoUXzAepf1/oqO5eAb8J
HoxoE5U3QOyQKPlE51JQy4XGiO+zeynGFUbn4K3x9LTUE79iYKy8n9x0Br04B3Cq8D2n7+GxEmIy
VfKSyS8Kge+O4KHRg6yp0MzEfF6yOuraC/mE+Pdf/LhnT6XUI/CekBzuN82w61jfq88IIVWkPZop
dStbjVmM+2msaNSYCcnAqJrOy+qAGxvBs6pIDDzfAB+ze8OA06Or8AAWO55inA32HYLJQoparOsx
OeCBC9pfAwIuvVbrtshp3OdCBmecZ8xFMDsqqPXgCvJrVaEKQ7T3UkD65JezAhcbvuvU6UAL9FMI
EsdZ0gmutK7YwpQzcg0livpzKgFcrVXfu0Zd784KD6BIYZLlrzpNavDokD4V+Hpo0LFWkwlRm3bT
1KOCQk9hLL1jZOl/31aiKAKYbsCtXwRL70ghR/G+UfBfl8y8qWWGR2t7C3Ce4miqL93N4UD0mF+t
ch130PIOCsqNq66YSIM2Uaj1+ZgJJgzmBjg+J7RVDKxGglSDJ45vMkSZ+g43h9nEIIJBkUzG7ptb
GrnIqRaODTUJ7WbFp02YN4Zm0VEV9T7L3F011Lo3mphnN/aBDRF9j8AXIoETWTFbrr++s3ioqmiH
teIK21w7QAO/AVAptbon/v5Geo59J2N+Ncnpqaj1VD7pYnmfi2a061D3+u8boZRFOjHClzeFOuXz
YhdBRnYPllBRDUDQjkaYnRPZpeQuHO9R0zEEdOngWgRzqbgrutPRZij+dPvEZKi9A3t6oUUzOpj+
o2oAZAzUTj9gGC80IXMxRIZGICPOR3ySfXZ5egRYXx1jNFaQIQdHpaG+yzyh4ffwbOlgWN4qm1q+
pyZMjZrNEhJewjvgK1Io0WOBOo4OTxC4BdSH5770g29glWROu1Wr+WA8iULT4q2gYgjlJdU4tv6t
yj0KMlvFM1Bgtio6sq+jfVqn1j3d7KHlbQ4JSJ9amDWUUuCp7YLjCrK/gyXMslgxcGjurtM8dAH+
OuTt2aNEQ8tnZsiE40D5k5FJq2vjsP2QnkWpZqKa0ScybbFTq8xE1CndqjPHloOBeUKtwIAg32zq
1OAeWLM0HAb4snogRLSPk7fJPnaPkVhszxFqWx3mV20IIcfvpL4ATzmiealYcx3Wf9H717UTLMJy
zYJ9Tjmggt0AOlE+3kIX4hO75b8PSfWsGCUaPVN1WQj6ZTgdtPanZeADW1xISh+qWjaFu8TZrfLe
1iiRjLp1jp9wu34TeCVmWBEvZe44bN6+QT/20GDqdr4aAOR4qnnPmJW1DnMe1OvzTvH7+OYldKRW
5BW/oRZNFW/zlr1OaEzWIvXa+VR8l1E0HN8YAiAw5pXGqnEV/NrFhoPboqa7Zaz9Hz3A+m5D6uRY
8qxRXaO2ObEIfpD6ljKV1J7ekYOIBgW1CVaYezyK2gUje7UgpX3u6lbTynxHCRACyvzgqznDg7pT
bD41nL/vViSk4mRGAmXVxguWKlYRkIumalFZF2j4q0859QGtzFkXb8oEGOpJvApc5A8aVvEX42sZ
2dpA8qp8V4On+ZuBkHjSqmamzGtk3XwmDx57Fa+UilT4TUdC0IexBFWCzGIJoO2maUd0TKaeAl/b
idOkngxZVSCGTqu/+B0JKrLTtfHH8YVVsKjhc8MH+rtQzpWM1kSOu9KEGvthEC0Aq+IEs/kw4ZU1
RCfAe7hu3bwfMwSrSrl7iGEhZQ2Vy1rg5YhB7HQhCD1IGiyk57eeMQThNetmJxee+MRDDZc7Hk6a
nmVNjDxxDeAPFJpN5YbqD5oe92aV62Occ9zVswskKK97hkwP7RpJW+oJpsGEGIdoJ9gm9OpOaaOb
s8eQo7sF87e3eruK9DK25TkD6mSnrhWML+Y6fngnzUTw9QZaKgu3u3NhBs5BVgq7GSld10Kx7BaU
ULLdmVEH5Jh8fEHJ4udPTScMrQnNiiT1dwCGfarBkfVwq1ZVLup7+Av65PUcTKGj1XSQjCn5nQgJ
XsCMxlQZzNjejDXGIbWWaNrAmff25MlMSYNVH04WjrhtbFATVD5o33RLTa5deJhZ6A8zHJY3Uwfi
O6lG8JXpAMLD9SzIXU7tNXQNTRCl9FwLSAbCavvfN7aQSiCynYCCqY0Hxz8OBlIoIZThqCgeTmGF
Xg4VyPWXp9DumSnd98TaLYqqgPK/rS3RE70Pxgmx1Z3LXBdIFtTrDnrR+IcELNeFGpgHxfu0luTh
000ofUs8lyMSnHRPqI2qjbYkI5efIJhnUxJxxu6ggUODhMDf0FGQQyimAEtntHVEzE/kJeGNUs5q
OoiPXaS/Nd0A6oGDDncKk650usw2lPoR6LMsgo2SCAY5FYMRg4j+Hbls+HCPGfC0cUhUbFkgwTX5
YeCbcM7pB6NV6FngX4aZ3liYZxak3BgFk8lkm0CDB2LAt3jj3McBiHymzC2QOfYqwZzHkPDhYQJH
cBOQpp1gYO/Di+TMu2QnlZNrB8RwgeCHDvwi9PXusnifTigdaZk7VaMLsWDhCLqOSqsmLrtBbU3u
VBxBk66d4OlXFGSNk/coBncgn39Vrtpyx51/U5b4V141xn/tAd2UjDq+5Mxd0aZpATs7k2OV/zQm
iX03P3ghLj3B/NshVPZJvhYWwHBu1VahGSfx++bzho6eA6ywfdH7HRJlf7OdaTfRTCy80HnYhmuF
0g6V8UopUTt/zIXjHCEgr0HnpEpi2iyo+KePG/FJJme0N26bQ6Qt07KRjowU8NshRxiMgCLbWlOP
/IoV+Ezz+pn8k5+kM1fvyZPqL4RQSqeElYZr9lF7O6BG1N2AXlqZE7HJUCUNv5vR4qEzkniSiKE2
P8c/lZcpEj3YfZwpbnXZ0KbOhBwjX611sT2tINc/Zmj7XSILQNNMcd6/hnSBLTEfo4joYuFVPpFd
wXIsH333HVhXzqAA4j3j5x18g8crCEh6TPefApXShJ93UJPGnX7jLSresyJ9FY2mhM6m6QAIhvRd
Ybx+qwNUqmG+AqJcwLq6ENDqOF5/wgu729sIsYk3N8eiFXEF9lnnopyVuDEXB7t9q3HNmkMuq7/8
AL5OOcPOuwAS6gSz0bfzNFSZqE84WRjF+MtxL+QCztIDGQ0gINPl6zOnTAghI1h70Y7+n03Hqdqb
R2g8areDv3QUJvtztLUUZv5uFgYMA73BLatnHMUYRChp+wUT2w+WwDQVNLv9mAFgRIFWGOImHL+r
y3RO8wET51HhAevvUypTWAgpBzgzKBoEgxtQN+vhBQqUN8kOsRCqYHnDAT7RbFwNNCNzlzrquNf2
PurOCQDJ08kanoCuCuvsHvgnG3RWdEIm4ZeimlGkNpmD6mV7M0QxTWv6rDpXA6axrQSGQjuIw1pj
txLMciRrOv5o2GTZSojFhzFFFfDgxe7Lfv9nklcqLpwlmJMAIY5JgNk7LF9Wti2RtJ+BGkGhMdHy
ADKPgCJelShHQedP5pJN5P0ZMzJxlIfroyilR93KgY78E5CB9z4MuGDLXFuDWoP00olvNioqrHYy
11Fts42/8BUmNSgCxSbSGt31A/MlTWHqGEyYGo1bjzcp7aD/L65a5KVmUn1/LuOtgYBra/HqMzx6
35LsjvG2C7yGOyyFM4Kd7wZyOqPL88EqXmQx56Ulnarad1s/yMNscH10lmPZu6D7Ece252mwSe6y
jL1dLSuE9freX6uA9Gj8T0fV5rmi/yABjanv9u1FH/peUv7hjNYvPuCSqRNPPZJwPd5jAe64JPeR
E5XE545kReDvBNG+5iE6LXBCzlaHhVsK7n7Ni8ZgSUXcBlpwgORU+WyNcmYB4Cu1YmPy+EzA2g4U
XOA72VusA+Zgff0bnmJnDHYhrP6PxRWi+OfbkyPFUgn0pv5Sq3A+0z2VKNBH6bLXABxGzTzdikVZ
8oBr2cWKdSNykK8bVJhL5VggFLCrYnrPDjKtRBfFGOmTvSR/UIpJzzvusr9caPJckw+tITn/z1q7
EYOstfHLRrT1X1CveiB9YddtUZbuBGsfPaUedVM+pvRtBjKEQaU4Pwhl1ywMbpB/xaFjun4MQkA9
XyhDElXRLzCTki+yfwNU7NFv0aLqZohZMCVIQs/MAzT2dOyRU2NUdNQVX8z7yIvQC4Z5T2pUBoZ1
X789xwrEiOjSqYMrYf2V5Ubdfb0CQtGFyplXcNlyFC+kdhULbj2WS/zLQ61U+Z62Umk24Bl3mK9z
65kfW6pyQX3XyEzv7P2XGsE7RL4AptbfnktT0p9hnEMoYznTSyZeBHfKPRnbe82dOTSbTCtUyOvs
NMdZOs4YQNlQUYH1eB2nOimC9zdlL7w7QRKTsrepw4u5Wo66pT4nQq0andJmT5A2aKehzd5Bj/fa
g8Vo+mbvMBVuwT5NwHXV2P65dUFPhryIszEG8SwvTu910W8aSqrD0u4EOWSa/37ve1KXSicba4l8
IHf26Xr6ZzlhoX8ovzDlP8jUa86dLNa4/w2yWz4MrR7a24JWO2jAAJic2EASKYSeQch7m6KFwHBT
PasKmcPYrlI/qBtX2gI+CbNKnmG/7Rlt1YB2aFKak1bE58gGcV1ArInWf/K/fOm3L/SqRUu4z67t
gh0Ppr6b82AQ/K0ck8b7R0NJnC95ZD6i/C96Mgtw3IEKvTdn08kzRt4A/xMs2g1JIWpv6HkZZ0P1
X2WRqGtRTtfuiYY3j2Kzii8Z6LjlUuut9c4gvMd4gbmu8ddpTzopjuTfavgx99mLt6F7l73bS4Gs
fVbRDOx4DwHjCafzTWLM0ddtzxOgV6EUYSjanu7YXFWlxNHt4+7THkx4HlFICO1OhX4p69x2FfEJ
65BZAUGg2x3zd7B0txQx+hyxnR1EcU7FpFerSRtqkLLdb3N/SypVymaAz3XCkyqUCGGxNsmBSGC9
RPw5/zoYT+r+H/M6Kbmi2YmsPyYYogvWeRXSLaxf8rM1TLleaobSJC7R+4rZNvoaR9BX892vsSwD
zQIdPzxPEsPpPoi45qnqk9WcVT1BRAJBIOxaqeWEtwK09cBmnK0wi+O4uphCGrIl4KCyyN8kkvYu
HNfWkqnPP0WcMMMxq5ZSJu1k3OZeNwSLVL5P8Eu4FnOyl2SOtVcU+ikSTQrXC3uGHHDmNDt7uSGo
qNA5AqLk85iMFNwffW48XGN6N0/9Orr/xynwnukQl+9AyRgDspDtTFrOpu0pYPLodGPja05W9XDU
JfUhDScSl6jcaXBtY6hlUwu1q9oEcxC6dBSqDrArkMUCOezh6Vp545zQeNpPm9sHXUzA7NIsaem3
0N80ir5ry+4CkcWhRoIuHElrZYGb+YKZVuC3RoCvktA3H1xLKaUYpweJ2YvRML/18f/QD2aVnmNG
Td76rK//zJlTSNH2/uVFfRWUEaW1RxVfKmc1u8jfZKQdLrthW7gmAhb+ObxnluuxGYd24TD4osbq
2H2k45MrKsELNBeitq7YFVFHYYPWHxGVZ9oLhXKlLP0VeRbk9v5H0UP8XBzZhB3jBKydR04DhMWW
zkCl5KQ35raKcaCajXmC1+jVIbUKZJwxOV+Ox7ZHdO0YsJzM0A4+zfhgEoQRG2grDhT3B1q+3REl
VmANTEl9q/EJ2yN7nH50ifvtKfLVUcVeldzrBTKjTdDBlqFhxHVdYsPua9RvHqAkxbN2lwVg9Jsf
C4ee46Xl/mN5kcBeFMJDVI9cO+XzU5v+dI6DChGl27q1XD1peGorJY0YCjwOTNliqXDoYPgNHtNv
EfkBUF3F6fi/k3KXKigZmoeOZD5mSETiVGJNuRDa0+zWOw8h0P45jsWFCcBM1x3OwJ78eS0a9Bof
wJF8q0i+kjTHSgzBwsCRfW/jLtatTU6H7RaGNvxY9i1Pg8PXJJkKZanxVtZBTBi++DamJGwgIUuZ
WW5ECwfTD+w9cRyL2ckN0veZ7/Slk5mgoclocfJJwXkk8zHoqElrK39jBY5cWJ3ZrIggMMQ/vlTK
+ze9djKvXjDfM0PX7/+Nq+JT5937HBrOvq1kzikDjyJcjzGi2bxuQB8LOUFbx3WYHy8wpOUhU68T
4ZkAaAPZtWU8kB/o/9jh5YuooF6KkeTbsJwnZAclegy4JnZ9c3UH2OnbJpliQFuA0wrNfWYxGALg
+JCrsF6rsAcPbfzlMllT+dLsOzONET2uecG2/zrOaIs7JRA5RhD/lIYTXbL7FX1LgxxGyaXsHa2k
2qiuGlTK7c7UK2N2R7e2uT/yy/mTFNW5JWAPrElmMlbdyomtQOlOudaxscqXaAN3ktt90J9U/uO5
Sv11+N30o8p7KzPoEiZ3s7pb0qW4kF18V7nYQfTpMD6ZwylMOeCmRZc+7SynM1w0rl+53m7RhKa0
dwFnhTAxKIOlD7agFB3zogY9quD8XsXPqDekKfd8gEgBMf2Ewtgs6BrUwAn2W4JzR6sIehKB1Pvz
R5nB1t5YdwVAz6gGiLAgv3n7UiJYph8oeBdFTmZOU6iv/QsVwf8MN8QbUzSmC2NA6PITAhjTWLF1
Sy/MlekLgVpe1SWVXGeGjv3PX9DoTCGF+J4EBn57bG7vlpNCHGGQz0Kr5xf1ImBnwmgdSXxvKssT
SfKPY6YJZauKX40YhWftga6M5sqyiXcoav+vt4YFipNGf/xgszuXEuCQAGkOQdBBLI9pjp1Sm1OQ
C1HTUjH8auM83ffvvg/lrHl4VriUv+GezPhXPtG3W4is7XvU5DZE8a2JOvdHGUX/6IToQINJxsrP
9iZ59sRw/b24SjrowDEztO47bjromcurHOGSotXYm+7ea1iKec6kcRT1xHvYDkdyRYVPtHm/dner
Xi/eOUtevGouvJ5XHej1ubJCkUlb8Mr1vbRa80lIbSl86lCBYJkL4OrQHzgMJa/sKG3G4DCTTqXG
4EWIx9NR65C6oY3yz8A+lsQdU85ChAaQok/I4vY6VRMeziSRGjeHYmgJywNspel2iQCQ7stmhyGg
z5JWZI9nqXLMqyogmDnhOgCeHebDwI5964tDsc/6jxLAbKqFOP2WQ/7yzS49pHJs0L97PbHuaztB
VZMcEeC2x7cdBQI2vPPZCMv62B+xKKpYPG0xCTF4E2mJJ/5GDN4Lf4r1moiNHZD3a6/a2yajrxie
e4iQ8izk/ZZMPlP97rfFSZ1BfOr3sS3XpZekyMdut6OCT5fWdct3l0XjImiyCtS6A1dupfVr7htu
OxAMZ8vCNhWqUHsx4O398079lb2PTJfiDpQt9qjH4Atdjj/QZJ4Toi4jzA3CrU50vLiHsrdwo3xS
Eo08OLjYUPU+ELDv8m1PD2Ic8Dyvs7nV+lyg6dwFWRuCFr9dsSafb+penFpa3c7CHg4FmDlOLdTj
qemyFOYlRXzBEXGruqwUD4HzbWSZcHNKDl+jUrkaxFGuxr5wlV2+ffq7xU3RHCR+LVR01Oq5TGka
7Jn5TQjYKh0MSRw2lMxYiMtzf/tbJ4miwd9lhvNx8qK9axPaB3Q20HC6F/6KhJFdiDWS5j9vMDWl
pJkIZFUffLVhTIoL8QTfg7/p5uJcGszLyceTvn/HWumaYd5Uz7PuuzdqOljD7OWBjl6Z8S1vKO7g
wNisJwRCUT1kkTgSWEe+b5RPqzmdbeTWNocaFvzR6JM2Z6zbNAdAjUZfM9ti4YQegDJNffugWU02
xlG4Xz1UibaMK6Qhdal+tpT1vfknBYnpo0P2zctEMSduBbQl+rKRIyqrWrRWVMdMW8o/L6qmy+Iu
oC6aDXQ99Unc6APe8c8b0/RdMhxNw3+d1qhELzNdWIM4ubsFuwfw0xKzJxPLGkGOip8ajNRH15Bh
Z+3rHpzvXvrAXOo9815/v6I5MWXua6znHe39lT25Hx6mdkcHxTFUm/7AWKAHQ6O4lJkOL3LoX8Ae
lczVSvnqm5ovJpxdqf6BD1G+1VuHod97oBzoZZRoG2YgNFA20LpaET47a3Un+x/Pm5VWvXiiMhiP
sWgQUx/UjLXatjCKFXtv/R9qczOIX0IyEDyak+b88wWsdyt9kIWU4i3aUznyDo6srL0HBIHhC5+K
Lj8GJX6sqS3WAUuZVJRl4ix6Q80jGWJl9KthT3B3g+qozdDR61MDEIl7SgZbxG3R9f2nNpBoX12K
hbwXjis/cxbnf+RDxTDTt7rfDi74Sb4MZtBrGJGLmsvDAa3aMs0Ai9YoLdNZAIth4KX1BbGE+oGA
v7tdn3HhXUAhr8wJNScd1MVgme0t9hIGpnZx9WBBofjQ7Bg3vgbTRHo4AWWlwbHBHHCwVBQ2+Axp
TY5WNZ32sxpmvQTrdAoNmXd1DK+aZO8K6uOKAYamllFJvGqjN8Qd//Cp3brbUIyHaKT3AQrxwo//
4RtziIosPceWRhANhERoNN9Le3kVxCl/TmE28HML6fYinTh2/mUkVItzhAaBXeIKy2/QYoGEVldE
fyDYGIfFNVM3QGm7SIJGWJ2ETHVHp/NnRQ1NfEG2gXyZoJGY2V293UEupiygBeUocgzRNPpSee+3
AY5nHyrptBEvJngODJRt6Pp7e096vTGRfl5faleAF9ok5cC9hjIAsnk6fkIyEO2DW1cGUmEpf3Ek
Qs0f/pvRGXntchkIrJ8TJAugNMTs6019wb0jjPqjR20A3DTTJPfYtNB2bjBDqSpbqhd0vbv50L+K
D97G9X/1C/QsEc+p6SY0FuYWf1TdTbd5unS1/jwDSfnV5wEVNbn+hXbI2wQQJgNsSTBlCiwxPETl
VtyjPqXkheNeaFkJ3GcHtCOuvbJt1IaTMoJMwciC4Z4kNa51/Q4Ng/Hw5n4W0VEpFwy1Qob2Fw+z
2bO4ujH/PWltPNQOUuLtstCpO3aK4V37ifiWIrVr0eqMz19W64Z17QZPhAd7zi/mGP/ZO9JOO8+v
IL1dvActgtVVLQKaYNo0SXNfUm93r2BIW3n9orBcKBs73onEQryd6juVEexf/pk0q6OF4UByNDwl
/HhEj0xHNh4kkS1rZFXaIfjp3b6iDpxo+ZWrvRmMS6NV1LOoN9ob4PPZvDos6dTjOITJe+PoRvS4
4RM/rGZcHI6AMDWYLsAzDDU1VMcOGmzPQTQdlH4VGj944qVGcBlkPgkO+FCOu4nd2G61hEi3zSPa
uppRVh6dX1ShEOTqooZoQcFj0OIpfOoLCSX0hczPR70G3/ta98DU0oPo4I+xFGlPLi35F9sa3cK3
KKrk7KToKCcp2yTSzZgTS92mg+ZR/UdJcXakw7s4lRO/gGBA4jq4lcrC7VTOJCedq4A0aSvzW3bs
TbTA4kX7SuH3NNPoIj7luuvQ+RWMPAvoBM3VDmCmWQh15WOTdo2S0OrXTw4uaMnKouPTHRYQoJ8f
hLbEkmUWd6gkYvbK6/Q8XhBs5zP5BsW9arrOZRF77+DMJ0ZujFq+H5INqwKF4ETKH48s2FrPZJcC
mQbJ2e3/fBQq+rZ/sgXanP1jtET9Q4D04hb4qq2AnJzpGu4TmeKrXyD5Zi83mvvHf8oOKIAtXQ8W
2M8tGk/1ZDv6atNRjmTQg13oX3ED7aSatfMkqIYCte513w6A8GdYm44E76h7uPWFX5adWsq9GXy2
nLRlIzTRnafQW2b71Uy6t/NxMQBaSlYINUMtnsIjbhngRmLYhNE7oUheAf3ci2+NdOkhguRrXEnX
E2QAgNY3Vwn34I4Q/S38v8ha/EoJBYKVdaY8w06Zn1W4oM25ci45hz+6+t11sZ75cWnvJrdWv/JE
akVTzWzV8sJPtD+12FHy+f68UBXbAE4m0CXJ+4BY9Jrol2C04O2OnQFGVFy8yhtOAAnclgwt5A7j
xQ5kulLejrrPNJt3n3lpQiye8pWUw6Ezr1NJHq80v9m7E9f6DsulY15oC8ZvJ1pSk4OQyYtJAo+1
O22HNfACv59xCJZ5t5Ar7ZyjX/62FUtf33UHK3NbNBuQfgFnNS1Fr1L870kO0/wYEvo8OPyxAfQW
neP79DJUSNR4iCVwV9B2hI07jAcTYgoYcRExP+DxEcMWWCMQX/ufnn5QJ2Mm7yaNi2kblyRPxg4U
JyBLdlsMyDXeEHqNFN0AKhQkiqhYWEyZwMBQOqAnKHKFUym5UMaPJH2in2K9dzYLyMl0uD8N1Jvg
2z/EdrAi17hGYuyQviaFd0PVpo7oCWVipUcqO+bVrKBhX4WVs5iQHKGfh1AcZ2KUigdEnC9q8388
OsN9EfqwcPWzWINO5csVrW/Mm+eQZCDbJNGC8nf8FzdAdbEBSLpZuJjn1WRAa8oPv71M93MKrZPF
rjwReg+h+6Nv34Gma9K2caDIJowDgQHgFeJCsY2jY4uBmFhjH6mH1Bnp3lTY7AiRnXS9cbsAxQ4q
tDGpDEYrNJ9ZCTNPqdyH793HGTcSTwAkXeiSbDFDLkb3bQkifHr4FWfC6aapkkVbXrxKGfH1K+rX
IkmTJqe9+d0akczC8FHw/VyWKDvbKgMqiFYOYM0q/AVouzZRfQkt6Ov7qKfZg6FnLVKsTmgZI4EQ
MPGAM5ByOrbJS47mrQUGbdy9YtsWlT5m9X86X5SSi05D1vd9nCMlIhahdkJ+iF5JC7/jcrDh0AlL
qXtcbVkejzJhMeZeO+CZCFaBBrDUkoZZuQmYGOghpXYJk/Vx8bSfX6ARgRLBK6wlE+vP1Hm4cIHL
c3etMUpxsb66rMA2LogLHsbPmMDm8Tt/vz/wwCduTSshi8rny4zSkr/DhYZf10vzl36Im1dP4Uz5
b4oqiVKxSj47jR99XwBUkf6sE3TN3ZjLUtQGK898AF9BSRHTaS8H/N9NoVMlVNyBAZVl4ePUDaqb
bL37xcuEVvudD+/azOlGQ8xNxnt6OPEBaBexC+aKvrpTMtOUtiV6hm9N3Vbpq5eueCkogqtt+qQQ
RBmO3Eew3AfR8rj1fzKCVAN7t03Tyw0VSJcG2CCb/2yBj6JOuYqOEIeI+yvmDh1Ae/jN5g/xzpT0
Bn/NE7rqDh3Oy8n6aV2ZQIhANDZId+ybhYpaUH9bzoEFt9tZt9URNNagjOPlIDZfKyRY3Aatd9zr
ojwBc+sSuquPdcC7Y/ZD/iVhfsceyz6lBvZgq4Z8CfFghLzDDOT5W7WIk6DS5ZP10bOt5U4+zr1b
s07JDB3q8WGVUrXqq9qdsxLg4Ty2QjImpbgCaQTISOudSzvWnUpoGyT4EGWZV5f1cRUmO/HvcXNQ
JUAYaaTC/JXOG33yv8AHx0KR3niS0sK2xQq0X6d5nBPgWz7+t38tEgX1VR4d6mcqVk0S5YP3vCh1
7bRsVXjf7Ez/RaFIfBSQqZFNKklrBYwet6IhB6b6QFNSRRDbInOAOQevHNEzcw89vzx3pciZO0AN
DXn4YsXyhJV9UFPvTJWkgmHu7H3hS1kG72DZkDIlqpz5DJNSeWDm5yKMna18ey5GQANghFLM5Xvj
zXXba8Mj7dpwEFiqV4VD9NwD0PbJvgZ3zzEatJ6s4uwcCXjQ7EboNQjufauWtpE/ROhrCWRQpy+A
lEcyViLJJuAK1e8zs5klwuUOWlWPSPMr2W0XNxRli2TD7OaCR1E+S5MeOjKkptDVuotBVGJ0Zin8
LOpDCCOzXINz0AvzzAH0vinMK3b8cw/gsI6LdLqTuVXjSdZFTW7BWAOlq5mL3/SDKqv7y/K1ZbJF
yIRIeCkjM+uXoNGeJjuPS1UUKbRTWO7484Dppti7xo9PuTvlENR4ajpE/0TGP6quKJZsdmMZ0UnX
PWNcgfPiQiURLyfpkcaXLnXEesNWXZUSJ3nvz+Fcsj+xdgjqKKXyIVBdDVwER/ua/C7nwXAfbjIJ
8K6o4twKIkX+iTcMIOJmZyYBSQ3F/ygK211OzKByWRUFwzl0rOySpscLeTXYNlTDUXN5yK4mLpoE
uIQtNO8gNb2X6mera+X2g25CTquPblsYCcgsV1bCkLhCWJLyo8kOSkX2EDn+pXVsfVueayu7Dxlr
bbIAwaBZMUCXetMOaX3Q++bEMtfP5VwFXk7s9FXrzh+/S6Sy2KeCzNGRDSuUH86HfQ+tIIJxar76
FpvVhh70W0XL0ZaOY0zsg6LVRGQS1tdKOUuObKSRA2gtIwxNHpcM4ZWDeIlBHjgKNQr5Gn0UF+wj
EynRLntjimmXkcnRZrpOHbruSzTsf2WSIKsO8NssuFIMQh9p/q5zYmE1/mgFfXYsPTJNbGoeIyqT
vVe04DKCKKSHk//FN5t+JWRa/Hc55fCL6hBvkIq2VjeeV7uKBj95UtDVozj2MqEPyKi6jK6yoeME
ucgVmapwyDQZTrsH189YwxE5EbZz8xYNbQU4cPmJGyN2xVweLkIl2PqbyIVfuJYaxrRJMvB5s9c4
FNgQnuRDT2UcZHuCbs4sm66OF3kqK/yzd55wmtwBJr83zsczRsXFLG+eH5WiSc6uItYysy/pMwqD
00vFxpHBC7zkGDuKk0Q6Hpdyf0fj28Ud5TtCU5aYWnBKNIqOoSUPGvmiU+6R2s7NpKjrttAdMvjJ
8YRPbsDtZUm95WyReWv1np85//Qg+Th0Tns3/s6Ve+7Q8o4+vHpicKbYffg5TrCChuY5fX4cnepq
4lHLLazO1fXq8xtosS/VO3rbJC2wbWB7YuNbOTw7qES/NybN+g5+9Ggggjp5kDiO/akOM6PGEscq
Um2hXzubl0X1PvDCT2xIDhKrCZGn/rH0QXiJr1IFD9/mgA/Ndgcy4qO82yKBeyFWXmCRvVBloSss
6/IZ7c/SfOxUxHaO6nOSCeCYlb6MbVTO44sBaWN1nLImkDHXbvzfVKX+PP5Wc9A8i08Afgt5kpt5
COGgZZ15K0+qrPJ0+4VB+P5Xow4alL87+SxtY4UUujohJdmcE5UsmU8A49uzEhG1l1gw+wvciTPf
kDGB1hqlUkwnj9ZWJqVx+Rx6dIKs1o+F0rF/ZtT4gHSJgQASaT2pn7FOmvSMDMw6moJVFMcEZLLE
tTKJ8Fs4/yGVtqBJIzCsk6q0iR7wT7AiwzDf44A41H9PrvSWTet+nb5gmu/eXCljYQ96K9VMkERo
JPNWtJ+FctibdkaqjD4O1zxXrZEXBYeGKTAJvSbTcM3y4Y+6V0RGyP//Cy/OylUBQ/e+2G1Vw/1q
O/MTSXm+0+2ltxOq5Q/8u6AGZoxGwiZ/WRRwRQvqiDv8meHF0svgMNuSNI6vweChgcipI2yFIB/N
kjRcsyAm+JV2Bzdmbue0KZjQpi+m327tkdAutUvOrtrK7DhkjVKsFI7wQtDSQY9J9cFQ0RE6VZbk
eq8R4OqOvUDoFocgUiZDdv0VUl7pSb/z1Z7U5CdxryL06E0ew8ppu93Lgs0MgdWXZR5GJ5GEqjom
ka74BrgoL9nrynCcMYrPFzat+DrPI7itRKiBtFVHz+eJ07WOutk1Jy85t7rJhnNgKwno96S1yxUv
S1qZhzRne7glIrjqrLdYwQrCvN692ISqbo4vsJYt+6N9BqHOV2XK+3WH+ejPb7UcnevwBdgdyjrq
ZskuPdfP1+vtD98FrHSET1dTT9aEifoRMoWdmkxwHfP8IPKB/wbjxa2ezGi4GLKNBd3j5P3lXgQ5
WDHjS+Sa0XyeU1X/Xweuqnh+zxaHU0+fW1HNNBfCq4Q49GpO5DEQwZwwYxkDWj55b2ZJAcb8X0BD
sDnL1WYFNn41KzkPqeyzC/JZdPtOS1+jtCQc9tpRiT9oumlMudIHQPtcrvZ+nIsGpRfsFA2ys4A4
TGD8oKzUg+xVsBxrMPjj3kD6MKmp0+5cnssp/XsnL5sKZBpAo+lkpodHcFcC21rVoYo/ZRZRV08O
ZmRmO2Rym7Wm3GDDIMjZgNj8/o7OxGZXziDMEci5DO1VqyqZg5rf9jNGzCkBkljrn/+81muq6UjG
JSnKbDBqhcrmfWZN/cEOGkoyn1oDymXafyXmIElljQ60szpU715o41OqtjkkTA4ZTFycQAtwgmk+
FufIN4nZNvtp+9GsnGLXVy+okaZIvOxYJz3t9RWe2YB6fyv0PhXolh49NfOdEYL82ne54sxmkbQk
zT0OKQVQE9HuQ5PeNGZ+G5rC8LFc6XvP48dDy9GLfoPzGQc+dYUzVW5u8t1C7BB/DGVkPru3pA8i
Pq8VoaSxfZugKaLU0krc4OIZAOY6wBRvnIMgJ22PKkCEb9iuR/WAvzVqcnChWqwzfGICXXARg78k
wgT/2ygmScBZpGWseKC+Xwk+W4W7Jf32Kug542XnU8Or+HFqDUhL1dNRjKrc2VZdvGW3OjdK1ymi
SbjsDsO5lu/GUnDdQurdNdyrxuUHgW/QwXoEH2LhPav6FoS7lyX7zZeJlSOeWtqQ4VftCxeaqicx
n7uujgS0dhvs0G03q0nhQveurFu4b5xAm1YMN5Uh4LX/4eSgirDtuRHcyfXMlQE/8fpKUzGmX6hX
+sUMMtRHX3NMnOzv0T9klj1qEQEi1g5cVp/7GfjDnDGwS11NHBhTufCn5Z0Ggya2vSBUT0vXKIjG
3Nev+v1t7gNBtsIkHbsITSkJQPtEigapSOUJmBvv+Y9PLUyK3+UE1P6RsVzrhtkPBU+jshkfAhW0
HsJ8/j8lrQs0DjS+ZssH0lV+meFWpo/uutOpMsLi5pj8pzJ2xu8OQs2og2CIA1qnvgBJzwfPQ2np
GjFLBJloUTMpZEQIc3sUji2cpGraUIE3okmNNNqBXkiGSF7/YeJdo1kqXi+1u7UA9jv80AzZA5fl
Bs00rBvDv3nlIA0gMQKstufUAkpPIUV2hxgoFX0y/iAej2waKwDSCeD+vFWVUnG90qJJ5F2Zqf+v
9vuZnQIB7FfN/oIROh1SqTFXywO/l19o3AQ7J203IMXTbAzcj7CoYGeIvPY8qC0l4Qukn+dOVxpm
bI9BjGEfQunC/lFhkqQflW9v4poCTPnMOmLlwRQ0/Afu6BWDglETmDoSmqKPhi8EqsIr/Lg+b/C5
5WfpG0Ofp6AjRFApUTfhZB+YnadzAomwZ6zCqH6v+OWibficgQ7/kcq0jwmvksKN+WNg2zPQ4tfI
k1q79hmeuP8L2NvCiFixpHwAcqJXzcWX0i13e71hOom5TTmjwpvgTrv0w/gDZY7HWACKYNh2hPZ1
j+SMy19+IiAuXiP08vDwdpILCYbwOIHNXENxDAG3OmIu04u5kjZifl8oeM8mS0TvrkAEbhyv5Jcr
G4tIaKyqJFfIX6AOIAsbiuxA/gTbwoN21na9CxFC7g5qTW7m3dQ52csjNWbQ8tbRVx0r1fNC2rhh
7bcv/wUj06/5ZeP5WvOOVSInU/+g50TblHXSLSkJlTp34T3dupGR+uYIifYzCSIcdt4NujA/YVOt
G6qcBb3WA82kMr4iM0kt01Bma7V8LIJP7pIwCphT3Js4m3v3ms/DmNjULLY0F/oEVRSm+W0UjH2/
uxdqsmAj44M/Y6uDO0AbtEybZKpTyyv0NX5JOfXgfr+M+1F+MnveSNiGUGCAzoa0VdwhalbLTXQB
HD0gdFJwCJ+stKJWifh3/mxVRdaRgIm8qrW0r1bCEiXcCVR7892u4bu08TrUZObYCwQt6PzE9Y8W
3nRg2rOsAfOIm3HVyawj+Wwb4dtZ9FSwgGCOfmwhlDVX8BWwm4ofR28tvHTx21XlYlvf7mknPV7Y
mRhDK9W0+rcKYKxL77OmaCIg45drFqOKRtQMnyqjXRiBIHGyARlTeLbM6xctcYVhBorATIKKspTe
1MM1vbbcxZKgP/9/OTBH3tN8FgUpnNuvE2HdHOO7/Doj4ule+fkXLhCAMrtXBGey05zWlypEzwBY
Hi/QsqP9xBqxYe6Ebx222GdriyPPlXLaUPB+pdNGxNmS/SDQSbwO/LBgqKEeX4H5lULSSk0lB4fm
RQEUxcj5DPtmN+iUFAMh41uFZ07R+gmxZ0OvzvMWCaAHpPBcKbXJgQWaV2YxMpeOjJpZWo2B7DhP
PFdGi4UiIPyoiF49Zc2b9mvxfMf2YMyDySWsosjIWM2CQ/9Woe8n8g6iGDI1DCx3Nt1/sAoUW1/S
5WL/waLHXOHdgcuuhsOdgDOfd48B3gO1KdthLON6eEF9lxPG9KaQR2Xs9GBJBTznYKI37gLh2qmy
ggMJvShTudwQdFrNlLDK52D9+qUXM7llaeXLzN54XVDMNuqG8NXgL+ZI/oPy+QpINwoaS3jmLevg
StlllT0yp/F6KizMvQi9JEhVIbTwgl2gTtC+rxZu/a0HR+IorRomPR/kYHa48xJmqavbUuf4TT/J
PT18u5+q0LCTvp+aP0qpc92ZTb7nIm0fitovcL74USiG9vNC6geZctkjGu+EpnXndFIdEXumuSBr
CGwvG0fUl+IloUvS3dSQqeOeGQn2czv2hwyPHkoXFp1hSTx2KHyWbF6XSFEiGHCSf6DuokyFxmxO
NVEa5s4K1GKycq7hS3jaLzok08fP+KCvqUO1eIeug7p7qDvQombeCQ3LBfVyql7/QytvnHhEzi4E
WSu8m9+VLMZ+Zkln6JCrylgXdGS6fP0qNh5tEWsQ0Us8Mk3Iv+FFpS04SiyzJ/UhJ+8jpJlWuNdr
vIL0+Dvylq1avfJ241UA1gyusgEf4R08v30oPsaCE9Sqe2166UzTu9jCrPOdI5ybX3iqB4TASFdQ
bq4v9ihybPskMoYkB8ElWkS0TtEsTkpSpBJWDFVku/ArRmSjqp5vyESd362Gdh1Oc7YULi01+xqe
z0wHisptUdK2mhyUIa7u4E3AV8TLFPsGvyyg6cN9fpzFA+z0Q3sNmQOg9rhtgXIQHYTgh2gFNSMM
o7vtw6k7r5HvijOXksCPNMGgJLllU2rGnWM98+ggHSJD10hns8VGxsxK2bcF1qI82exuE9lIdIVY
LrTARjmOqf81dndQSXs8AwEpIigfzpLDlwKEENDJ8h0i5r+4DcN655Hr8XnaKnR2Ge6irMHaiGkZ
PYSBt4TL9SvYIZQ7OtpfvRv8gq66EADHluD5/C+l4mC4e7P3CvoLzO9jTyETifYOMutWiBUIlkoC
4a9M4pNh/NVsI3+aw2kiAnt/H8IEvL57BhJWb/AbCYmwp3/lFWDVB/cvj+OypsA7c+JnVrVFI34u
sSNOUwdRJxhtU2LGKx+oQKKVD783cBgHzHLDQCb0bXfWM5p31CN/MeSs4NauIScww2wK57SyR/W0
QH7Rs/hd9OSNCOQsl3qJjVH0QmwUL9tLKstTp2TMQ8vPZmfM5EwXVWBzOa0kOiVOR5fVTJXAKKoy
yF0NTpiecP7NY8Di8QlDg4deWkTVFbPaGOkW9Vut/nvZaJwokLzQH9wz8Rh+p6/2xwVp2PmtodZ0
m/cB2z6hK9ThW0C7DJ8iON+RcKwJOttsAhYq1hjl8zdeOKoxcKVbN5MiimRLnZBOP7Yw79l5khhQ
/NLjQRUuQ+EyLQ00N7gITqbjCwYrDwp78KbC36Eym5L473Gwt5fpdzytxXRgFdchzY6vOqaOeTUj
SCTOh8kWbYP/cBDKMgqt+XLGdgys1RFhfmekaXCaFZiHqsvGkcr+bDJZ0Q9tCD4wLWoWU4Mk1Trg
pMNB2zOfSUY00XkB0aiDdzwhHHtCgWg5Wt9fMqgXVgSJqm0VSK/cdR/GDWnU0EL+IYCTwWuSEst9
+Qs6ERqCusYO6t6qjna7spnQwRgwS84gSuNT5MysWyBevfXReIJywexS6BeQj84hpyyYC+KSDHP8
yKwth9QCSgYU/bsStLr/eDTVSkHg/oBnguWY2ToXoCRFN7cGE9ZNPxRqV9FZxcuRdwKi5snXiXcH
UGmUU+RCws/ll2/f+/Q5DsazREoFcpZQKk8wT7Aap9MT29WfyjX2huNMleD4YnxYPHwzrZTf/FE1
wlsI4DpK7DPqUOEbzt/9Q1hF2WifLYAihf0zfMzOSQ7mV+WDFj1J9U1Ok0ihcVXXcTcZeJgyCPJX
+PMMV1/lXF/XcSpnskFAuvAk7ed5U5PpJKtnpL2UjmGNto9T6NbeXXdOmlz55CzS4r/SIvREC5we
gMiwyUGOBezah3N+x9Ez5bgl00b1Qi1Ohq7eijTq4tqxMbVghojsAZrP04NLH+hOI1gTsUTE/lkz
X1m6CEpRLwLasVasykscsGtrvYSa7zKfkwwe97702Mi8QOd/ZveSYlYFpfl/8sRlqmUMWhuKwEpR
VyfVVotTdyKeb5960FJp4th/cGpiuMnypJ2NrfZUiYXdnOTtS+k7Mfn8KQbhmV3GmPoCYZL/ob8r
RX86IE4iux+Uv6MbFcrV9Yqg9rcjDdzDrE2Q899f63cGIVtq4PMTToAsHoqcoJ2HTJ6M62o579iS
UVrvQBe6YF5gGEsYcD1PSOpaHZw/kkvlAEqnUSmmjfHNuErq6jV52Zlh3pQB9ur2nltgMB0XTWZU
NBcRgam6TAPRKmamrJsRMDiIvjoCKovsDfyv59b36If0eH+yohXslqOy2Ciy6KuttRgWX6mJJirs
KVFV9k9CGFg6bD3W8Nf0TzI5WIt4+PlvS8C8nojS8/xMWr/LihqOA8CmLouJ4xft83uUT5Keq38z
iEFGjgtlkMFuvwYqjcnezoBLQ/83cM23Ki0miyQE038krH1I4eCxU0BY3YTH5ryoh2AJ8aCaf2iU
fU/KQQrZSIj3ArabYymd8/gri79s4qK8W5kL4nZo8Y6t3lw3XQONcavaWFsUTeXPGUt7CeVGDISq
oz3f/QJvQcVEmpisI7IsH0PDft04mVp24DrFPfDhOyhNCYTB5ZPCJzzYuFcRHkFHvNap9k+S+E09
4oql/R561rnYMFxjQrYtENg0CFbMeXO+++ZM0pHn+cfxmYvm+YsZ8TnoZeNunfUHa27pWNfBe6c7
uoHIivv3GG3M+qy9YGJFhyZCK2lZDDSgaT69YDY9AGynujXiFCubiNdx1g1GICQMN/uPF2e8NQVP
9ykLy0MsRj5gwbkLyXKC0iVReunfJ1QaHC5aD0jXKsvuNPsapS3yNFJgDZANOt/ijx911ma3GeLw
1KYE58QLD8EwYV1os4Oin/iJek76KWgm1CqNuJlEPFvsQPVFBtEfxvI4NyrLBtX0bJwQq2QtwUFh
+1Gjc0WINrrla0KpLwd9yBsD0GPGLrwXj7thhiGJQ54r3vRPobTERx1eoK/LMGdZEj3jNQRLU/0q
RIANIgKziFfcLQRaA1pr793TF9ASrgbkxeaHOQIsIFJxb2l9rcDzwU8TNCwbqFPMI4o4lXIuJwgV
idiQAKvQkHgSc4e3P6Squfbkfh2tvTod86IfESNo3XLYWYc+R7v2gWBQTW7fhHNVrlcwrNwJUQWF
XhxxFM67CTKwyGkjPTYUynPsx/Ajvh7W2d8nO7WpTvzuTE6HD31Xg9t5St7GZXXYXdvbpj9MYllv
ZuNP/gfGlIDD8XCIONbT07OP/WB2kFvRstmSjExPAv0DEOy3s4ylr9QOXeN4mLNOhvKIiqsYxOS7
vSPrGvuzwySD3wkBOKz7Q4HimY1m9YV0Gt9+eehjwQ5hX/Hwf3wAI2VnHr3qCfbcI8wPhN0yj8YV
WR7GJenfpIz8xpSeAJeuhkD2+gmkgWJ6nxb3An1qZQxTkpstqN8DXMtxefZ1lITsJzIrcG16p2i8
aJoZqSx2KsrrI9LoY1VMBB5dr6y9Oa6/yRUme1t3qUT5C/atpxkOF8hnvXP3PRdTGBA4Rv2RwYT4
16+UXaSAM8oFM40td68j8NUHvthu/uPgKz1geWJy7nGwQK9NUOfTI/rbZMF35tfXIRY6VYneWfdg
sOISmeVfBc9fo6ypGkN33KZY1R8c1f0IWFBx5F42SHcb68GBIZ94xCusXddo7nuQU8mShWJek2cl
aMBl8C8kAI1BKfzUsXLGOkbV50WuXNd5gG5M4nbV05EgGgvWaXEew96/W5I5PxN0iSzzYghRSR5q
LfwJ0y8jQ2df48it413mATuwPx5u2YUASH9GW101EGoSbEdD1KRXhundHz1mHqM8HLQeXRpf94kV
A6SMPvHVjep1n++04718GKlqer6Fw2OR7CNg+ghqi7okF7zIReSHFslRmtPCK8pfdowngkw48RF5
eQ+YTB2ZcPAlb1bVs+Wr1sETc8MUpy+eQhno5YXxVemIatoGSLLx+2s+cXNfZSnFhEMIb+4xHCFu
gZJqTM0BRgZ4DQnBL3VL8tUFU7fkS0RgKiL5mTNxX0kkOvfDNkqqiPW8/Yxguu5HLaT2XCNKyMlp
+26V6q+CWgVTqKU0dLyOG0/POXFt6Q+EJaogeVidAaCdLH4J7Cl0oohdFbqq9l5WVye0iYMm4oiG
qDMvgLFUnAiWJJdy8wggyS0FpUfv2nly7YkkyW8Rm8ia3LksCWyUEtFeMekluJ7H6rM0PZcad8Fj
sHUZr5+bfoidMFdyyy8oQqe0LcmKd6kiBpqT1FU6j3kPCxJgPO60XVKREiUcd65Hsn3AqVOIyFCb
QI/Wx5DEVMDSHaBhtlwVQVSv2ljT/A65njCPzuuSMErdczmepGyM0GOz+GWaIqX83N4zRzaI8uBZ
HCEcd/MnFdRHIvoiX/Y9+hG7w+XEPjpeZ7TlMFLxmMoKbqItbAwKW1sGoG/GyUH9BjRAOiXq6u1q
Kd8Oln2HKpxYevYkvUlt7Zu8gbWOZQhxXF8L++csvfGGzimxKs38suF2tDfxKiFt8OiYYFR2cSha
mud6AfH/hkCzKHLTtpKkg+BfX2BgSd6jwr5POSWNEv0+ywXjQMbuCXfphZ4DwRsDmyUnYBTwi0Dn
01Y1aYqH4GNbyjJ7fAwFj8WmoVSCxdxB/oMQ7aK4eMm3Y255LWwm4ui+dt/aJO9ZhE/n3xzhUENt
RnvlADFyOe6/S5JfN/NGxMvdFtnd6vjr+JuCMEySlMwoXwL0RDFM9jTKSJs67mPeqPCoq+VcY3BY
QG4S1PZy9ToVweFC7Od8wzH2gR7zshFrWmPqaFFk+574BsZfx5ZNCFsLWjcMLxGfMb06yzV93BSe
mf23x3Vn/bc1YHPcZOV49Bv0wm7BrkDih3K5EZh1DZO0b413I+SUNOvea44ARITBfEbnobgvNuLR
WiO0AVn7ipBzeeCsl0weAS9JO+JmnM+Zctq7E2Vzna+e/dgJNn48LwrO2BKlKUGNog9tHH/oQb5L
VnN43VvaS7ScswfFOiQ/gaEOS0ZZlA8rhoPUUZpNWFNnubKH28EoNhANHCm6EBz7UbKXYR7+yTWp
HuGep3XCzWtoXrlCIdXylTmP/T6BcRWYUlmrEV5ME/34Y39pT9AJLWjv0lbOvy+XexNSxYdto8PO
8h8xBnd3JB8apQl8mWhkeTI6li01+R5+P/cPTRhoBHYjfmhYZC9B3SHPQTN1AO+DSukoAlQQnu4H
7xIoNgp6D7vUtJaDSBMi+8+PDeuwgxy36I4GRgGzV1W/Yoyegqrzs8JcFJLzOwkZUY/y+b6s4I17
buA91C6eENH8kzEnn05XCQmUyOxjxTZF/0bP/CQq8dAEWUcoeum7EqB/m24QhBc8QeFbs1vX7uX4
5QgsohMYc7EZC65La4cpomOCZPNl/2dJRedyispgEDp23KLdm8LWEGuYFtrfKEnFaPUmWDeOPK4F
AquXzkEH7bCzMp7QbItZw8zV6SZ+4dtCF1WnMDGmgPQ2dhSQG/3QNwhGar8PfRrVmZjEjCLNJDIN
/P8DoWOWOYrlRCuotYjO1cW1vJqenhzt/80nBRD9M1NtIEzJnTx2Fib/svJqklbIn3J3ITYllw6J
ECMiW1SDdTpBMq7BPrOpCn297USfWQMaDNbUvemAbFGOfk7B7eqnj6018ZqyKZ+fjTMw1bKXO6Zh
nNbOQyprXtptJi6Ksx26IbeXGNJj1cpJyNumoKLxBIA7idgKdcGMi+ExFoYAyv4tKSSr9TcDmQUg
ffe09B1NrjXW9uCV/1s0Q4JzyiPQQtK5kkvx8IAtmh4wx4QTj8yG/Sh4zTREIisZd5YLgcnpLFTW
bZdgbZF8NTv5/ss707jd24jdEG4NIhkRrhHoxyBm6MaHrYjIQyWb41ymyDmSu5XBa/foZo739jp0
TBK4dxc/hAvqCKJPNtQ0LaGyCP7OxzWF1UgeN3FTRRzK33hoQgphJnzsVkaklkDauAf8/hqk0NX5
MrY7AWTOB9acNrks52ZNVEhmcmDflbzz6uC6XGbwq8MeozkVsM1TuiirvJJaJXLMhpwePtFQEelD
iTJUnt98OQk+89Vp7hmQmbGOTk65ms4l3cpmnn5ZPSOAbVt2dw/eLltKJ087atvH19UTIg/eBAuk
KjUKbigdh3g9CBqRsl0Hmi5gB+RUbMRLCm9JHAEF4eeoC5UQcx6H21c/1ulisw2FBvxn6Nq2uL0W
FSzspwSH7yv9JTIUhYMPMqWdLhqiMTvtGUXBAXpxVk4F7e2GYEQhW7JU33qhDNihFVcxGVo8lgat
64ylJMEnb/BKjkrS+P47Mwcwy4sHWt480nV910fMjKaO4tUZbKf8uc1R+2t/xOXM4y3oXPakNk9j
bAbmvmquGodnaj3LeO1aECh1sTwyLAHH3SHA84x7WTUwU7F1X1EuDnkWOeyTvu8WLIySdo6ospIM
795/wb0cKMui79+jil6r5F4U70dveAOelpTqfwI378dDGHhxjbNU0d9PaWkDstL7SK6OL9D+IzYd
8eVjBSUIL/q/rMI/hC7sL4631k18waTPbhftV4fMUXhyq5BVe5pgyqfXRDP/BHmXT8IMVXPZYUe3
r8QRPCMluaeVWn7kBdyAANmrGfOS0WBlWeJh7CFfcjVb9KcIqwR3tfsYBGAUvx6wjoPQfLyC7646
NaUiEw78JhSe1vsaZ0XiO9AayhJkSbqqgkhUOqc4WyaL3PUkDqNtsxTRKU2E2fXf3Jbk8aRBPvOp
hGGi8LSxmwW7s7IzvTm5UdgoenpX7YZmp4x9h01lBTmt5w1rKqUfokdL5P+awlycusb7jVAb3o+a
DMi/wu+/DDFLbStLeGj1Svy93go7MmkWJZrAJuZivUyxe6gTY8OjjqwazsxBY1c5FmfAzZTA61hd
C3M6sd4hP4zvvbNzGJ2qc6wPKxhNaSCLd++B0Qgepk5wboT2Bozo8cpch//5YFIOz3TM/wcs+BIR
dxPo27EdFH2Smocg4Mi8WSgZig6pNvkpVjMWcemJi4PO/8tuxn+DsKVsXBUBfB5CwBPfSvqxV4xW
oqplZn00sT5QuzRhYxyZyzVh0W5hWW58wXZm15In2krT8R2F2xqmd8B+iCtEntPwHeWqEAmgIxKw
aV4HHXRqr0bmGh+Y/wFgo6YSgdWpf/Ge66crXahj9zHBjNnOPNdWHf5D69l3IZWHEfeTrMKdBSZ7
fYHd+MyMV//bCZ252QuemrlWk7IrO2/KrLkWZqZSzwXAY7tHBpbpi1Ee5VS0xYAAIGilFt79EMNu
iDuBriAxLAvpPCmsh4imGJesAsu3dQOgaT8II3k57qTQQx1UxFqy5+kMK29bSaMqwapHuxigy9Y0
ezZXmSlG0FfawfySMazzcltFafOmGDZDC3ACZ8tIi1f/O+29n3Q2+Bwp1rtM/Gd+FuXqMELUl07o
KB0SJxALQd7H20EvvoR2H3JD+YgiLNzliJOwYJI0C7v91152WaN+OpmXA/kikV1P9SdlKwLWkPkG
LpwEEB7tbNIhkhYVm6HdsgnA7h0r82B7bGg72Esr4o+a91TyiYJf/bhlXg0qSLW729q0tP0L60Ol
BbHy2O/+Wt0n4m23DmlyYwVz6nwCgZW2c7qOotIFydtbqLT1go919YtB+qxlgxFzNBAAjxd84v+5
wtc5VbzjDN7KQDXyxb/pCgoJKNSTzbDr+x18Krty0oKySxZOa580MdisEizh/i+BueeCmxc0TyMp
/iqfrThxG8ereLSpPk9iGYR5wNbj1x3X7kGlPuKk+3lpCTwqUy7dGF3XyWNBedRzuMPOfZrLp9ct
3k+AZIGduSsx+71aUAV4xV1IsiWuFz5rvRnnQ9+j1bUEWB1yycUQQvkvBrvdiQ6mHBl9dfv0cov5
5ue95ylzkq706Bjyq0rB0UJUL0AdExkM0FTb44DzMrHrovXC10LA+GPkwQ33ORQZQdjyIGuouHRv
8bEQ24B2qsgcoNF6aPF9MNH5gYhKmzpNXeW5o1r1ox6q63ih1VIBP1S5tAKCZDoUDrVpJ9bvPn9u
YK4faL/LqHsQzhpN9dOpiIgdmPFmEwBdc+L5a5fbEgPGgzrRqq5hrZjL8zkYo/QDdf9+XPCt+mk7
wKuIU+wdNARd1OPYE/6q72tT+GxSlCNHVMgq8MFsQCX1Ld8RlPfTvTuTZ6UKIukwyuU9Zl0OcAsJ
cOtTGxDiPFKN2kIffDli5az9nufhLnXmc0u6x8BoWE6rW07flzEUogjyWPjKzz6ONl/2hKjkmXZT
XRkd4msSjZlt/Ix9T/UK2m/BEZf47PGCBNB8Jxv6ucAI847OyaUKX69AynFHJxlUYXjAkuXO9nLx
iI4hvJ0OLiUu6dldwK/6LAaVhsBSQv6nQgJorNVHj4A8gvzHrizJAM1bOOkgVySs37xkWd4kdo3d
2k6MUO4ZxPNuKbI8u9P/SupIUbCTK4B0gJj+dMkScuYd93O/ZhglMKZzrnQ9sTzmg87vioz6qfQm
zQkQAVoqUWCbV72nyScM343QfPliZ6L6bvvc9p2IKsEPqrkydgPkB6UFvXlZElR0fOyIc3XFvbr+
1txsR3md2obZV8zFTFME7gLBtb5R9MZoXiEH0J3+kCRAHXWl3BplWsL4jB8gdTvv/aPcHAJbwOC2
DxwIN59xbwvcv5E7QDldMVQVW3hSm7t1FFS2Arz+ge+yA0eRoRg4uHw75muIYBOLB2wGw27AN8jj
KN7vrce6/Ha4Dav8OUygDcns6Uxc3bmeaB1jzQNjdD8wh9pY1q9bL0mRKkYYwR5jbzdM5QsF5/YS
eplVdIRDm4+7zsVGR6dZdXJNAe6WM4At+mOd/FhKALAd94BZnVUL/Z7ZtDe2tmYA3MDpHvt5RILj
IFBugdHdmbOsWuW4LUqLLkbqmbUj4WmGLWDFqkHESwzqJ/jGLYStAioXBaJd7VhekuPUMkQQLt/K
CZgLABWhYykJJAlrT6beGjSYxaiyqr4+vKUIeY7PtpdvvoziqRON5zlXg+wDIhZ8lEKVLNFwSyBZ
fH1w/XyalTUl5ccxmeSq4leqUSRandeJFpfA78bk6LZXIGTioJkt4ZJsyR8dhiw/3+Bk3e5Vs/lO
D7kx0Jy4BYCdUMAjQmoGkg/ZeJ9fJCV4UQ0DFCQHPyqYynsj6I3vvTIjIpLO1QeAtZx7pDhveTph
euq7DryXVItNb4fVgl/lT77TS7/+SlywX+C0jYE5qV7T8LKPqvjB+t/klTzhmApBxiyjGK+1f/KS
ASZNIK0U3xG5+zC54tQXtcJtKaT7SITVJ3aV+Qh2EbE6Tcb6YEVW9VpZngmv2W5U9Z2mH++Fo0vh
PI26tyNTI/L+rtvWUahWa6baeZEZJ++orLfmXUnSPMh9SIOiXM5vIEVx9fd3EvPyBN/qq4kbvoht
ZxjEEfnwwnenCEtPxsXD3s84jsDdRoS9hCcxxw6wWdYee6EMwo4eiD/Pn52XzcHop9BkoXDfVFy1
ARSlZX+VJbBTsdfcQaNEmvIeSjtsshtq7khcwRXj8PYfYUsY0ILIkneVGfJZWWjcwAl/ymVEzrMc
Noa81e5C6gz3itttrrMr+RSqsuTmv24IIJuWnAvAjrq7wVyGQ++PRs9VW6ZKMdKNCrYvcYeUd0Zv
Y8wP2XaHixwunnq1ntCXjwLZnD4FSGBhd/CYkyvbHvJYn+9oYxBf1by9DeVzU21HwR3g1Ej465Sr
l/pynleXapIlUCwmf61QGU04FMMMIFa7+U/QpNquQEebvALMSblLVvrWv/0LwgYQbcvs7zx9v8lg
unnktpXfgN8UNCsOwtlOCkF9tkGFIHLE3sxu9EPeolm7YPk55wOuBkks0o8CCX5BaxVGc6D4Tx6j
Adt2+fV+DVtgcpufcJGrD+zAIZBUg1dbMR5KxYQcb6AEM+Vvn+sCrFwFDMuuKqI1LoBpZiaEV9Ak
CKO+Bh1QIoSpU732R3ATGlFshBdYeqcMVlR1xfWhtvv1rOkAJClOYUUfXKJAJ2/CM4OwFyPVGiUm
DUivJ9HWy4fjoIghdw3wWCo5TEvM3qixYCBcuNVNSPJf4zoEjvAuaZ9gCTDds9INB8hQM9/PtZFM
Xrz8RvyCyafMkUGVxVlqqmEzojUr7S6Wj39lIFHy2toAEGfryqSHurv+NHn09rFVZZfHZATKIKGd
UVzUOr52emSmvlqUe/Fj1pirn5lO/HEqf76jYgYeEvO+o2XJ5HD8kuW6by6Q9LdLPVsjdugRecGK
IDAG+F5Hn1J2AckxUk4Oz3XNPbX5y70cYkzMV6C9a+78is4PoWAid4PwQGf85sDgHT+q1jJx7DGR
OuSvxN5ruQlXuQilAxcXQ59Fd4GQh/o6pmnSXGIIJkWtV66RvWNLR8PCBYXgluS08km0VFoN9gI8
6GpW+APqeqDzXARMhePVZpRBZmn0xOtRNByeLmWszCDwXRuIJF3TGFyx5P17uh5oVxmQ07aguEYN
cakgc+9KcwRWan6lA8a7Fjy+jgGeJoIPtwJHzE0tn/lyXMLB/3loxwNANA9LJ9KGvmdzkMgOZd6v
IDas8gk0KQhQHgLAsMEO/dLevMRsn4lztgt7hvPhcrSqes4AtpV+npzTFEe/t0jcrowdfj4SXZ0p
0LFQuUdfI2owAfvra0i/RTJ2OHQ9HQ0mrvjJKA4r0WNVWWYe8m4eVn+0LVjk9E8XATa4LzKP/B99
XAv5CqoaWiWTvRc2kvz6a86VHKJTaNz4psHt9z/OJOTx22Yq4kX2KK5/vgJs4bwr4Q0ClMNNnVOY
AtFAGfSUCA4ChVak5dYGmr2UwRLxvdhCo9Q27MA9gpWXo5z5cxa56xGTCSdI6wpWww4Gia+llcnX
pctDESRLA6PbhREaNKjgwEErrutx6HSdH77D3gUAGyEEeqAhWXrAUUR2h7689xIh2soEBAlrhy6R
9M5FzEAf6mISpIomx26c0kevTebC6yuB4maD9EIoNdzmF/AYJP6BjfxlDyjIxNCiRmsvwtKnY420
Nf1/SAe4IC4nSMamQhj670xTYh48I06dD7017HWwmd7uijxMDn2ggK2bOJolfKjBv2gjMJuPAbow
0IpgJF7/Mq0vQ+5FF/8I8L+PLpUW28O78LgtG2qNCAw9TDaE9LfEf+D5JmIjFB6r43+4F+4AyI5O
msnf0jzzeAJ2UrI0eBCxJiIlLfcQfYajUy/nwl4h3Ceow3Vr/twRj2x3XFiYIl0tNaHlytf8qUT/
YghG94Rlvq1MavVgAlrtckLo2JWMkBa6npIMDw2NDHWPvOkSGExG3vUagOnZQt2Zl52yniN00yHI
8pJk8XLywwPpeSuij9FdQDwduAu8g2M3lI0XR3Wp3uYeDkAJumUzV5lcKtRt0amzqD0T6HB49S6f
pEeSi1jJT3AZ0YUt0N8T20LWx/khHGvk+Y+/ql/ZzV8256sJJqOAePJPE4e7VSnFKA1GWHCGj18k
HXptZMIB5boF+tVp11ojDofRM95V7nenUVXJjbUaEhaRON0TLc97ekH0GYjEK1/q1IpkXjM1m/RQ
GkCQmCfIYlFdhI2XgOxHvOeuQ20yekqzSiEvps5q64pvQeh8+2elLlPruD74Jc04gv8FpiaVKlC+
OhCniOpDnRFjNx8cB9yqntyXdN8+LG3p7Qc/cQIIjRQH9rCLStZadvgWCYz9+uki5jrScw2t2iLV
we76IwGHB2AN59zttQhDicLr5lYuleOmeiqTKgCgQ0hq1UD6JdsdlqcHLVQhbhDf+s1BKlfYbzUo
lEkxxcQTjRqfZY1EKiJOnVUhcGg7tQqaxsjaubE4hf5+b2ZVMRVkWkxhOh4KJZ+jiFGedGRwL/Uw
3L8zqSY0bAzY/vyBvG5tcPdb6+NzqX7yCty875GfMDb68+jLhyuQwA4f+g3yYHL8tmkQaimeG8Gl
TVGXa+aDjWbOKDFGiZ0LcAeZoQnlXm+JStbOCA2JDEwY4IMLLl5uXCUUCqTYTmLPUHeNIKrJQ7O7
KoJC+h65TlpLXTatFYEBRXrR2b6MUSf9+qHaDzeHvcFQH8B9eMo1sMwhvxuoQxL/DIHYkn3o91Ji
lmngcmndLXPfiLcTZwCMDwOuWUj5PBX3FLTi46aPZL9rb1os3rdl9X+PLOf2JRmUprNgO7wdDgTA
3vfnuyP/AaFZAt1I971T5cSWAKXFsWaVRuzxlATMUKM6gcfSjWouwLDUI1B5Htc6TdT0r/HbePH1
O3RV7xZa22L7w5khP0dJXjIqQ9lZNiwsAaKUUzWy1AsK9IVi7DteP2xniZzm9NH4QEYracHZQ0HB
rZ5i0Ef5+kV65mjnVUibBLtdKWpdpcp8UR0x0FmLvz088jNkHLbZS0lG07Tnx0daafHTGCa6w0lB
P+ougQN3PmLFHGFCwz9WFppgfD1PFk70zTfhBqxAq7PGDd654KN60aBVSQ80Dt/IpLHJBPvxsNON
3VkCfvlMASo0OnMxez2ly4PmAYxzUbglffLCbJW7Fuj/YDHGRtcSI/SVThOvI6NXjM8UeJqKxo3v
0f1fBTvbI+M1Q1xZvL81bjCEN+hA4F6tC+B2l3MezT+afBtX4eyQDtC4BmBu/W2lXRBU/OR5z5ZK
tmjzUHdNrLmJdmT/iUYnNnzNf4THK6XyKfG2RvmLPOrHNawyaLCbqnoeJTKtLGtfi73xJgfxhTM2
9G+JMyEPZsN0CPtoF/WcJtnrjgA3vxD3GFYWXiF5RIfrBUteo2XYbjKObCk9Yj64SUDq45vh560z
oK2M8jliXdxSeQKYPCJYkWn363ok5bQajolNqtaF4j012dGBRBq2nD+OJw678Mpc/5oHTUjCiT8O
AO1LjeSqDrN3EEmCOKpCRBVqqsnmq9l4Ew+afPHcmevrx3Pzutsacq3tMn4esgCL1/mgju2GbXGw
of9/wCn7l9dLMD+aOQP+A8yh3s4tPw7V4jq5Ig+kPG3nw7ScJ3F1hMCrcvbYfcFSJnhhxcLhsNFA
wXRrL4k8sg3OprJgPWXV3nvHUCsf6kdt/fTHHz0Em6p07VPT4t1u3Cqs2K3pbhxmRWf54Aiga2i3
TpgcIRdgI8wS6Dx7yqq5IorlbN+UPcWtQN0tem4ffG+89l2VoshQudDPW1K+Z5SZ+iR2gqQLY6F6
EQCR1ueG8kIlkii2Eeq1CmAcbh2phCAijtIq7h585SXx/LfeiVxKjilgCOe2f3lrkMJzaZr5XQAn
wVKhETX5pCpnQKSP1kwnAF08GA/KyXM5vOVcKVgRLoeWRwVBspwWLAaNrZ5Z34qxR5Z+8ksfWom3
3KE7cG803i+ilzXsC6pvxV9GPug2E4apO2iZQo7K0na3B2sVyK/sNGAXXAAjCBddWpYnz59wNdXe
xXJGEjPZRGAB8oNrEgE9SqCZjyg4IwEO0Ie1NH0o/H/vB4j3FpCRCGJ4wj/ScYtL4voxMx17MTOL
QA2ksMWJQhHtfT8A2N0xPv0xTn63i7X6+Qyk+NEaozNf0YS1a40HSTusnI/mnIioLEh3k8dsWuyl
qI8wyXsM3vB5mVID+BL4F2Q6VJuXWoLVMAzGjIFsFn4BUn67OhapsU4bvEhbU0yJJFt1KLfn22bc
7xfvlW0IrYVuD0sNHc2+QMZj5C+kFEeIImYn3ThhKEG3HV0ClOkOTSOj4Jcn1DpL9q6kH6DYBWoO
02w927yjUfTUQgRcY+u54W38yV+LvZNTq5XmXzHb5SYx6n4YeQNyRl/m2MqubW2JtdcZ4FAN9osw
Dgmnh92fZNar9d0uDwTeh40k0DlcLPD9YPbLAH8hN87X04dI2/9IBqcUu61dzYayrx33+VqMrU8L
vRNf9VlWeU6skjAphGvqZZ2a0riPsGiV2Ve1MSyzNZLasw4GgkZaoLLJWNe6g30gk6qcVHucDNay
6ycVuzfVJrN8HKCntAU1l64eKo+AUfFqf2KOOWa3sVjRA3+igYUyazcWTG9klKZRdHPCw+Y/mgWr
o9A6icR1Ebc6HtI4DadpyLd/vTH2qodfoNDUH6/myrJbIuE8kvCN+GiN8OI1hwED45DgZ0OSMXQh
ta7G6Ji5pDzuKt9Mzm+iWT5DtYsvlk9uzggOMcJQNauJLwfomvv3s/4JWqqSwdhiE6HpC5OSkJ4O
hUa56Ot/+bxOJKYv721arexVFkbflgPXORbx+OwHQd66S5gqWlBLb0vxHoleP8Bg023xg4uc4hXg
lfyY4rpXFHss7hyfLi3idC2DzZpcnQhK/E+wIAXMEDSZfM+zHlNIYxMMtAjAYLJr3Yt04g3tCGw1
FqZFh8NTpVZN2wXV2Uxn639dwk/lB/ryJmknieSfL3Upu3tmokPv8ELRQWLJmlFRZDnDvnMJw7ld
zvvjAo0xkEj2VBEPlg08FtaDYojJR37bZJ1UNoKbeiYdL+vjYhfslzSuP/jaQfGJ7q2aIxMGWY7Y
mdJfNiLX0x0onX+a58jc1TscridhQMI8zQknV+0uhEq+dNR+2si5dq0FSgsZX20IZqvyJ+bGtD7Q
+6YGowFLwFxk2Ns8MSv1C/y6e8rHMtezjrLOaS9XLM0ZoCA315TQsZhXjGwsrN+0slVMWYE/H8JY
lu1ec6xxoW2zuHhuosNnrn0rboKipKwvEkNoHlOPP6JH4MU4RclZeJneX91MivWlYaTALIFUu5es
YbsnKBk7YGHZjUizyREGYvMXOfAf2N28XqI+z32iQjzzjlGill/nw3X0bQ8vLStpzgHcLEz0XOBm
kF2fnrKW7uijtudYf6d2qZBn/JuNBDAfLRQU4FokBU42DOYh4s8hpQUDLygbAj9FMn1kmwPF3Xmx
KmxPIfHkeA/Wbokqq+RY59gy0Yyz1GSVLwg2UfdzwAwisXMB3UAHwFOJOS7/MmuSPw19XY4y3Z4d
RthVosLTuOqGiEeRa2iK9NTq8atVtBBvKQ6x4F06VcNk2M24uUYGTpaFOznBRzNHD6YlFKc88hGA
dcGOMACEOah5GVLACJDsXNdO3Nr1OinJU2vMPnuUyV4ZBhr2JmcE0T7HAGhWSrbTfdIWRsUW+d6S
AC9qgdTwe1JfTapx0Y55wjtueAcfYgQeQOrIDyScCUquJ1P0dC5Eoa8ik5O8PLuEQQyv4WpicHDi
/oQCiGVbcd0TuZwjt6rbASBg0NnMMZJkxy4piVZdZ1rmNur5mFgWhmEP7BxqAnqKeQXCv2ihbt1B
Mo4FMcFjFTDYd/8tlJHzEgI4NkBMHoGjMbq4QyvY5LfeKfKUEjf6SXWkKBYtfrhkfT2WppEBlgjm
X9K0AZDLqHtl2uDOZJbfYusuh08XBv13XwM8hFoaVvNkdDZ12vEYf1TwJWtqLT+YYyn+Q85WJr2T
JLfo9U9aaQ62foPwym5a9K2ktfwK6U98yqPGN97EKqXAmZ1F0XzF49hLk/6SIdnWmuy3gHOZsuLD
IbxsDDrWlDhkpm01Bn2zsc1V/GQbloiZ+L2UJ9FRZPoI4mq7ClrKuwqjDQ2ey01eToHxTN/bYGZN
7vPaS57/ewjVfc/fBW0UTdobv4k4/SqapMc0Coq1HFUa+cLevUVg5jPUOZJX7zDRXNfVD9/TrUUF
KxGeA5W7TD1WVYxnrbwkIV5G+829ip0CuDH4IvL+ehzi77UVzPvfwVgLVojfbawRnDL0kmIHTmMP
Ep1sHA3jLu6jUHARBkakoZ1oSa+y+chpTxSbH6b/s7kBWQCvfOZuOR1Gkrx5y7zbXmFEnl/s5v3V
hyDPK3ygk54Rsu/SKKMKFdgAoAH0qC+oIDrJNgGjJRPIVPubOmdczc45QWpchlcTT0fJs7rZ2VP/
pguY8s6xAbxrsdBX6gKUVM/4IBXac3toP3rkr9JFIvi5044Z8dPnT7J0LSTnrJLV4adq8bIEvm53
0aw+uBx1AaaL0Yi9k5VUpAECYw5zhduS6VvtmyGu0+1aNg29ijHilLpCzKym300QBIIIMaLBF+cX
cUCwcNswYw82DQwBa9yzght1MQvtMKCivMn6ImSwibw7cT6zjcRqU+VzZsMxNsxUmNDPWDqMvaYU
TgpccmagWXCNUnY6s3xd+rtrIw0+TWqm7xjQZ6aARtT22ONh577NwoFOWF5Q3kjQ9UEh6h0Rofbs
zAe0Qr8ZmP6H/vZqzXXI5TvhfkSDtwOe2HSStCGCj+srRdNKMxsSDer6hFVDHIrBYN7Gb/aqbIaE
h7SKbixTNhjM7dX5Oym2d6TGtSmPulvZaAIwxyjKFr6k8tLt/P8505pSXc2ceu1mafHgnyo6/yOj
/MkJDql9LqbSfSzuv5wv+VzcBK0Ssxr+gicyAVJyD63zajschFjqK+hv9nLr3c3MuamudNiIwzy1
FEOB9dBpPrFBLDrXhwPnnPRQsWBZZCp6AqZzCzngYjzbQ/SCkfzJqd7r3JaXEZn450H8/Ere//M1
1Hl61uJAgPp15vqdhfAFUIM8ifBr6SJiyng1nOgckO2PnScIpYP2Z14zi2UGpLq3qQPFXXTAF6V0
/UkGdwsw2mdvO3dbkMjt/fHDX4KibgK1I7PvIfxsBCww/xlNoBFlByrkyzgPOZCqteuMK2bGX6yg
r12apsIaRWyTgHpyLq8yq38Az7ACnkDYMBemO7tdlgj9Y7rlIJelIVlVEJQICpH9tbsYwSKqzR71
8HnIQSTQqHRG8pxYmKTPT0S8C4qaRgjYL6P5i+4n+IBj8ILViLm6QcFP4qWWobQRt7XFMWUrdOMq
W0+TJBhG4zRhvNPKtiHgxE5qPa/w7ngX2vCJm587E9SLsg1+pBo/VAWN5nGHbqCgtunrpQfL1+K/
c/46KWdHkhb9/rCdjOKCtkrW/kKar1NjwvIcfBw90N4b/Tt6SkQV/mkzbmECggfK/Bh4lhf6sPiB
tCN06T5tun2X3nlAm42x64hBRO5/sYnNfqXoRTZbFud+CczNLQl6Woj2lxsH9OQSp4aMU7vy9ahX
HD1v5MaZl5WclE4SyYMQadKpUNubXUJ0WJmhsJpOc1QHv9VPHhvij/uefVopRFllT2nt4GYrB/22
ATXjb/JgsDrhn4LznnEStdedWYMKXCGQbuDwKSBfFDUK4fq+sRrPp7dh95hysG49SL69HLkgcp2f
vZ+z99PRXtlkuB1+O/TT7i4M/vPOKBcPY16V3JK+1GgS6Yx8CAgWNwA95/QR3XhahJ/ArgsKPrxT
drxbc0k21p/2lp21l6umD/7SGbh5NmB+gXgy3/UPVW4VPxZ/WhgBaQBzkhaOTe7vL1u3ZZMoJ7AZ
k30HD8vbVhZJb4zGk6ep3F0KSxZ9uO+QQj60AMas0MT+Mdk+qpgyTDUdlwe40rLUxCRsSL/xy+y7
qKCkNE/HwZVhIepT9QVMPL4YCUCQwMEs/jvoeh83DR9cV96Z2xvC0LDbL4D7JVk9WSwLTXlItmWk
cZAqKvws4P8OV1W0o81iXI/JKt77DZ/rm2JiWmvc8D7AsphdTDt4GORqmbeFZvoHb85YFrn2rU66
tuSrOWXCL+kETTmjhnbtlEOOJ2udJNaEeqxTnIuv3E4F5qSE7Tn5PQac5FlntT3pSnRHvFP/5CHH
mrJqk1sk1J0W+sHjAVY6lCxlkDyZTR59V1La8iv7rY+pWAt74X203DQ/fG16D0aGMwt1DjHJRXsE
v42Wwm+MwNivrPAkylGQe9g5mxlIe8m4VPL6v++Dd7gPSiDxdu+lmMGBXDKczDccHDpautzCggiC
SMnDGOvhaaEClH8DemBWgD4zh9Uun2LJPHoTOYNOSvh3jkwnRR1ZWKmFBcVwliT+Bjz2O6iLpEbd
HeK9VBNUROyaGMOuJG93Pgy5YvPFj3fn1J93khH4L1vyyJo9JzxLHGuJkZ5hFdCGoHTjUc7AtuKS
i3UfLRGIT+iV4dDnkOZQGnsuL+jlM0wex6WMV0lQO40ETnIy44jiWtyC5kRLaFaOzTFF12Zh/vht
fF7UZMniHztsVcLiI7NkxByO2tZnE+7Qm/oTHPop6jVUkT+iOyRLQffftwMEr5hu8lg5q7yXnvIz
zF6cVex0EfNhvvMJRVLXJJsKPELi8X4YKNbd7JTtazRTNOv/AU+/DTGlrC5SQEQuVuJgGNcMcYuM
k6/5zu82i9pAlqN2TdUGJgT4aktACbfa3x5Jj+X3stKxa0fqye157HcRTicqSGZ7llHUTaEJbjMT
j3Nf3qqrEZeURUrQkTnQ5m0hzkT93DQ5xQJsY27KY4XhrppJM41xPEBOlSoVwpB5sxQnDNkRvVEj
KWusWY3afZlpzBY1U0ltEOTSuHjazcyE5ok4dETwgP5CnmCMd2Kjpya75c9q99NLyv5cC8fE/TAi
nvB6ByOD7GPqsjzGz217NlWD5mNqhmWf8T18H3SEYYBTh+QBEgj9hSVRBhr6768gxf3bHLDQiUN7
m9KyltP0czg7u4vwi7bd1KFo9qNnVI+CvCsYlkoCa2PWcNdtARdpCjsqEo/FOiCnxPCt1y5fTOCl
qI2kMSb5951s8jAd5wqHqGlAzYTw/cDJpkqdPkC9ojS4xSQAlVy6oSl2kWypezK0nIbp3XOM1P84
Nq3J7HJX4DVtGT+s0T/2nVdTluVsubGACH4FlADrLh3jUQ7Cbzl0gfCbvQxqtTZsQPkpqjdHBig5
iQ07RNcltzxJItx1jyZ1CJfjrkuK6xOlEawzvs2Uz660iNfp+qGCBBnVOoUC8S4uZEvCWjWbt3Pe
VNZMt/R9q7O48uRElRUAnD4p5IXNS15RJ5pg/Ss5Z8bD3yYUk8/sGNtNFypqljw8iZL60PWnEz8y
OIjk3qfLXq41wmSz+GyuZiDELihcLWnz66cRMc3pTWbmUd7p6QarKA5egOviHUM9M9XZtnxA4Uuh
KPDYp4FywB6fZRyCJn3tMer89Y1P8XuBevfGeCDT7CtBRgyaK7WO+M+m/rFEufj0yKBiirO/2BbV
ZIGPjfJUcg5dFIM0PDAP/R8C717rjNcIjByhmp7kzRs0f5jQODcKuZH1Nmj70xAEa7NIwx514qAd
z25oKk0PXVhcnJVJuEX4m0sfkbH2ljL4fVGX7tUJO6nfRtNgY3uHPCdGSULUV2PdW3WB0ObICnB8
EK4jr+Aw+nBJ4p8jZUutnZ75cNu0G8RQdQLzBjAejQ12GAewel3zs1wCLhsRt8iVBYnN/BS2myGx
w/wdrJoUnCzV/myL1qWDEhiD/d3O0AQtlvuBw02YAxQcsHs6KAF/FgO4Z/k5YtI2iLzkndWP+tGq
bnIYwRooPvE+wMOlyCNsT0owXzbq4ik7RpDFFRmOkbOqLzsbqk8u98VF86qVfgzrOSkEc/7QsGjn
JLMXoQ4xxRKFzwjYFiOpW8BjR4AjGgoswEkQmM//luBAblyIP0kjl4KHKaH74LzSqDFU9+Iyhx1z
DFxy/v01jixlhOqqaJMWOy1N7cR706PufPjIf1rVqq6AMqagB9akecHVdL1bH3Ezrdfy5MutxEiI
hn954CZpOZtWPA1WEfdXUReTRanHK58anObuJc1kX06fM1rAMYmT5fg4mAoQl9ydxsiZekJFJjIx
lRAEBMWNnXs/hEAY30U++i0PvDIoRECfsjAr5JOcXbgPwNnoxVs+JjHuE211QkaoWA34T//Xcb/9
HvjjrbfmRwlD7BtmJ354T3MGkcfhyDTqu+O/CywbpNEqhOoOOvOcug0IJ85KkDlcpJ5lPI5mNdMQ
DvC0cRtSjAQoVNbGekhcQvGt4mb3Q7vzGzIcjs9m1rE/AqVBWaXgYLVFHQt3G1jF7Riw+aDj+GQt
3HxtiNsuYhbwqudZjQIszTUmiu/yiNeg5jEiW6HM3qE7MbLLX28cFPBtx5XN5B2qgJqEOzg+ZblU
L4wEdaZZawpflbp7RSNtqusEvpG6lk0e0dcPyQAdtusXh6M4tpbEBp0QxAD5o3xf5uALOhspYVPW
0XcHK06A1nbd9R2xGiqAX9Mx+jVC9MTBgz3tuBx4EuOxEGGG8DhtwgAwWOPZHPjHPZGxQVA8DK2Q
0uS89elyKXgf6nkCE21uThInfVI+ZHIkKtVO2Oh3S4A8p4DoDVwLNdGCufuD13ymFT7mt3drEQ63
GFYiww0Rg8oc/MNC3AX09KRsSJPmZWtymzknHGatm0I2kKiIOYFlFRyESUvkiVsxUeMBq+Ck34Mc
ofTAoPSUUVk8xztGbfGvQvP5KNUB/uTiORcNjdx7yUHZHIBfSqMHf39fzefqnymwvDOuB7YObRIZ
U+6q6VdizTWD8lal277KXLaT+LVpkW6ISFYc1W04HPqk1uCov8WFT73SXPIE3gCeJJGQOisUUZKQ
NrcFFKA2l/lZSDwyansmQDdQ6VOVO6wy4Eme73yQJYExLqzfR3/OK5oaRxacGed1YC2jqx66Bfvi
t8bjfayDFaB0Zn9aFdw0nUSljgmCEJFKgBpLagD9/OdJZvhMyR/bVrh1ARG2JOrUNwVij9iDXVQr
AfuStTpRz3bkcvyAqDwduPrbn7oAqAcp+zUJDTDUnxORt+MLvZnLRl4WgnD5ppKAyIDlHvJ5k/h6
9shgxFSMdl2F3K0qJFkDNDN7YTIvnOu6jX1CPY07zC5oeQbo6NDTt++NC9DA0wPF0XF2qZCVK+ZG
twT/7eWy6+T8kYlu3wESoOuzLiYN77rHw9fzZqfaXFnnymH6A1zvdVe9I4fRWQQ62KhjDluyilkp
pdrZ912aFrvLvaliq7SC3vswSBVIjhmYkPRH6LUfyx3KTXhIU8mayZ083JnIGxugOE5a0oI4+2Rt
mDL7Ug9CcJrkeW/6OAnULWJ4yQUvZls9kZlr4UOg0JBuA95P1fF4DAwZR7ek1osyGZFIlo9x4wBu
EzE1iya65zuSARYNt9rPlGWR/iC5HYS/4ejucZEbVCGjTShHhXVLGNQy16GLshJpWA1WBdifuCs5
j7N7P7Z4ajgGX8vg6HAzuRh0jGxi9y7sWh5f9TVfJDLHDEN8+KrvmgzJOvtl7D1vQnQZLlJ6yCeP
EXL2uKWJjK2vVaoCmGoKDG1tnNhP2gxcBfyUleDGM4NKax5tIB548hsmHoOmXVQkGE68E7Z0Y4Ry
wwSSvE08rUjusyiEjOd73LwsNwFVznTnOGBFlID+LsrSOHqsoa0C7N1kNYEezMI/cXUe6sZEoElO
UGu4Pv2n7bLxwp7Xy3R9BFgLTrhdUwLdt/cqwfQ+/8eT0ZzHFVG1EKx9EZiTlP1ADPFLCUxTuSVj
4e5euzYJgBI5zn7AHxelWNFW8Nw4hCHh+H+gUYQbV7nQXD9JsEbFRgjO0FLZ07crMomMbQOdK9Ma
aDvlEOtzP91ofw9Or956M7PFG5TeJKw1uWIUl1G6fPgIPGqpTeGEfxGhcOd2Zw2KqeCge8ewL4q7
JgqtAfGOUJ3v0LgytbgW3DJzQT8hw/+y7qKfIxXz8P/OmD0y04fYhkCzVQh4el7f0RPBzgY0fyW3
D7AX7Rqp30CaR3zUZSk9281aQtoxQ0aFS+uSrJCEmQhgeGut6F4oW6uNoqrDiH1Ks0T7kODPcGmt
4TNvbfDD4E0Uv7Feoa0idJZB0NEI01AvsZMSDAwY0CrJToWcaupg5MbjVuMtD9Cfwrf86CQSZzpj
A3MfYuQ4qP1k5WCEThpxE3fSyz0QG5/2DeYg/S8DytErZ00xXiCvJqNbIO5QuGm7X1BqZ5QWyCIg
6GfM7pbgiSDbNZqU/Y7sU74i43XZUFg938lGNWfQmRP/QGKYLr4+qh64WE9BXFafOVBagRn4cMdO
l1cpC1G41W+d6ah4sFuiwpLrUaz35z6maoBTmpxL90XoSdN+9eXBI4uBNi5WnLCrOW7duJM7q/Hs
zx9RM0g/lyXykAWShQeoW8OM/gIa1UgKP25lD8v1nRqQP47argfVRZ5QnzcUrVUW+n/EDbIENS9Q
RzDlOBkBeW5pl3BeogcdMiNW+TuXAM5n8HJpngFiv97oautd1MK7/fwobekpDhlI1eQevyPrTzM8
npI7/cyS8K88npcpBhOGY4aHnBgN0GJzvKATrytdC6r0xz9A7nEC0r4DN+pyoKb0Nni0WxcD4LuT
KgEUMyTqndh3qxU/bZ/YbGA/22cH6eGJoalGzOGKyt1nrSQmoA9Ny9OCcUKd4Tg09vFSRNTgTZaQ
Lh6Q0Mk6Xq2MuNCzuDUy5J9vfDNRCdOQ033/fFm5Hp8Si9ZjTTR99BLQleXir64BKMGWf6z07HMX
GXp+mYncPNMILp6685cc6tQmSsmICBOZB9weyk8xcJJupzWuNkHMSdAwzUNLphznkAFQ+8ujhkwg
+hrVoFKNRlvqHmHg6NTV/rHGUtUd9PJygUJN56Q6f9BAEvG4k8x9CO8NR4U6cF2cEb1XtLOJCKm3
zbXbhpknrjJv1W7AGR68FuEYeK/GSrcXpuPSsWmBzN8M0slOSEZw/Ju4rir6H2i7TQea2fzrG7vp
zf34Qf9QwSVj5X5Ch2PMEEfzJsiIwvcmaJQc9J132g4nVSz5hWk7Sm6NWItMADKnIxXISkV3Ka02
/iaaXjSr8xUWHCOq1aKNqby5kpa2/zDn1sZlTXDGiWBpjZp7Z49EMmCtRuojUM0/FxjJ5+vxnFzc
rulL8lv6T6Ty9ySN1PahqO47Pox6qIwfStfooCxBIvJYk/TV8OuKljQWBrIMM/IKVePkbe1Cl8UX
1qjQyI6hwyHLypp3z4rCe8SLD2RSPwPCA3KIExDCTNbCe45Hzpu/DjgayBbHBr+wl5Ko0MGWvX3J
Fz/tuzNixmRtaZgRm1unyi6U0/WHr+cIRdp8E6uCHF7j+4/nUkHIuQC1SOsUsm/3PmKk5AeJ4lEM
mgPTbut+pLhuewFkiGBSmdREqVRJWWXiA4hR9qPz0rmNRiV2T9XL+0cFCsJbTllxlF/z+xHqInFb
2mVEzdkF0V6Jprnvc0tTabmlg3CBw1LhhEVZWvHd586DIQ9heJvJ1pl3koUe/h5rDVVMhVXBwGlF
5kkIMLKg16mf4lYHv6e5brjiedBHSFG7S6N/cYi3Tau4TAFZhHnN5uLpOFhqoLODjZEA7snjoqgC
640LaChG78qErjy169JXAC6HGdjt8G3rzt48z7shg9n871jW3TYr58+KIuirYaTWAMwSYWH89qMc
EijqTOEldKgkYm4fl+sXz2K59ZQKhQEOaw8xtUQWus/CuHgdiYpfIQlWW3WVKv7E2lyGNy2dZ4sO
8IakOlqUS6mECJAYsetH8TKo1q2rb3K8OsVYREgkzP0JQt7YEvNjLOQVN9RqwYj1of/fdGjPoFXm
g00vAMUhUndAqR0ADPVBjVwAZY+1H0c4xlEyGrtIqpxUHJLzmxQHONw9FdPYrc9IFEYwbWX3reVB
0DEXRnmTHtV1Lngsq5hrrzWaljoHdBt6AVAZUQFZjBcIE455p/m+7EinezrsfN/L+rYAUgV9ZTT/
x7vfBO6ZME0abM582X6Y+Q4VoyeCDKaTiGbAvXL6w5Te/eknAy/TKZiwSHyyPEM3nhknlc8B+ByT
cbCf5JvTIF+X30/p7/F+C7S8NuOon3J5lWrt+dzlLiOMRp34wevEaz8Km2G0HA5t9tK7Cb/utqb9
W9fWtOFB+ln5Ac93//etd4rqPLoFBwOX6fkj2fqVHl2CYe9FbdIPBltGJjUn4bB1Skx68/+Farm+
ADoWwiFqSn5eYgFtlxGUhTn1LqGXlQE+Rb8ZzacmXs4IXaDEAs7Wnp9IscEEwDqE4e8BELP+S1op
Qdjj4mPcv+UvyT/DmRxgTowfDDrsi7AGhDs8yGPg4wnvcD6Sxz3YTH7Wyb6PF0dxE+6gjShiO3VV
/+gCI1/Z2xZGAy93ia+7fNFp8qmWBsiAgWfe+rpyBer4Jw3umEBoROY1ER2cauBkpRc5fLUB0+Vk
+wk0ixV3+GwKQs7vi8Ru+pc/NEwgvOIw6D/V0+DY29Osztm0/0Pca+8LzWa5nBKWYiJrBWAGybfL
KaY0fxxeiXo31Y+OS26lLBBhDl+sTSy0JKYzYa/nWgayroM/Boj4R7KWpMt69jCCVOvjB3F1NZLU
trOFAYtt5zZgbmPD1FulbteQ47ThRTvnNGaLx3cQrHU1GMm0fZg2n/+ZkFUGHVQpS+HJ7SeQuXDM
V7LEnBN0rvfnPzktShVJ/5A71ISDrCuz2hBhS+h+BZ9NwS1u78Y7w3whz4l66MxWWEZvzc7zUfyV
pkVIvJMZ3We6Gyh7BzOoPZslJ7PuNEJJpvEvupFpxEkFSCC56bcGjbvWSuiBWWekUkX5CEqhsF5P
XUkffLlmKa6yP4LblCXQvq3fTdBaUqXipmu5Gi5ZR5F0zDZnhH7wHPWfhgX9MX4/CP7japQY8i86
MGd/IaUeAHEuHBqqLWl8zbXM8oo4DRLZzV1tkRIlesCa11TlU9iW5o10t/KBedIDeM401vB5JwcJ
jiywQJbHQ7Wxv7AtTfjWcqnZu4aSDiwChXVVA0vwNaXuQGzb+cXX044IalEShYcfPE9ryMpRXFtD
rRLoPSV7lkOdRR+4ikUiW4HEkgDjjqNxqkWLdUWaqMD0nI+6d1+Mn4/bJ0ZLTBOfP4lgvNh4uKwa
D69SJqR5v/W1Q7f61gCgyg27B3zkY4bPRlMnTNitDnwR9z15tsBWp0l70RYPI0Wn6cl6A3VXlhM0
KeNJ5xOTcIHjceylDomcXcyWLjyF42BlSMDNJrcaBSvlSq3rjmxAs/LJm7qulUDtW3U/d+tTkxLI
Gz5oKLVM2eH+WTAmiwvfNCaou5DK2mLlQqBZca7T/lzAqbBxtOWQytbK5Ud92KHUsH2J4B2Hj1y6
foAgQDTypnlAlBq9qFmQ4Um51y87+RYLHZsHf6Q8Z21yVGoUrJZ0rEOkLdBQfxZ6JiqHoSbVor7Q
8/TYlFdgPnmXE/krDh4a8rqnUok8N9xs6mPJuwQCBrFYNIDBhizFj/1ABQXXL4xUv9vKxBGMMnFH
Vk8ZD1NXeIx87tTrSkEWLIJwYHQbNp85u4ukg6bkQ5g8f7mL1Y56oQGCHo0F96j/TmoXxfDvE6sL
Wwl8YD2wnngD3LbBrYkKK6dpsXITJG2H4QClgoKgSTaK9Ggy2CkUoiyIm6UvQxDKqRwCdjyct+5D
eTbwuGtr6r3kjJkLFUVeqXAK56e+0JEz/uKY8mC+nhUBU1gWQ6XiaWGihO7jEWD4LXDFAubd8c2N
MzPK90pjp0bpFcbsuhnx+D073n5ig3/teuhEjwlB3vL5cfRxjOhDMj9ZkT3IXkI6CvByT4slTA1y
0FD8QzqgT5QL+lw+oDrZPMCvuQrKvIfHCpt386PzaquY14L4AFcivzzT6HNVFvr73btz60mlFPKx
51hSjdvhrkP090eL95/FqAleF9QllXQgwBTi27ztGlf7Ie3yxLiIJAE6qD0cGWo2nipjVOPgzKeh
9Qz1Lz6kbsCGmE1gMqhQqtV7bl9apX6KaCN8InGm2SKD0IRqFdBzwqXZwKlpzW/ecFgoDfyyfBJe
8L9J+wpLI6AnMvCa18P5iHtjTp9bMYd521xDenmKTmPEkSqyBGY7oNeopNzPEuj4CD4kbgMI3gU2
7n3vJzPifubbPCuk/2CjqNZ6q47j72VZjRclLZafLx0elWZX1UqJFZ7Nv/HA4jcjF0vIVjnxgN1/
uAVHSfIErgbrFEh7j3S6pyjT4w/VlYOP5oBZorvftB+4imtTbqKrXM/+r5+Hj1fQnBAxI0vC/nty
TAcZSpLx93CuXMiclTaHd3Mt4oodVtSBUMlogc+oUq35EdwRcJv6JnSm8Sugkrj39X8RSgVLAR5O
u0P8G9mMXxm4RV9/D7Q5T2oQw+pmktRJBz98k6/dJlrZ5yq9Xiv04vGMwTCrz3KPyYEYS/YtHzP9
piwkPgau0N+fUiFK4vOHOxpv+6OLxZ3VKFxuREkq1lb0Mx1LRmgtHpa9I0cu9uPSmtSw6xt5TXFx
dD9P3pCWxPb4XHPoIFS99IGnL7hAnt5FMuxjpK7Les2OZ04qQQQm9GNUT4r1DPcy+QcduoBrxnlX
+RxtrolLbIJsZF7cLsfRU8Q6gksPHK+MgXT/XQUkSAyLgcnZJ+oUe770EI9HpKq09Vb5cOQiqZ/N
HGm0GY5xHi2ciEpIxHIrBEUZ/viL4a484wNdslzDT+NuWN64uVmD41osFKQprWJh5SslFBNNOuMl
PCdmlSPGuyvkAXA8ykv99j57zrwEde/QFbU6FKEa72eOnjNLG8D3f8YtKyFrzy015ZHvnVt56sHV
M9Cb46+WByDnlRTRI/tCd628SaypAYMAR5VfRn+wSIO5znicebf51ive6h+qQoSzvZN8S0PB1QW6
7PBXdd7JLRKFd6guVlPR2rFvhEekjMI3RwWJ0iawL50jB8XJo5J5rDxIIhVgD/oxY5cP6pC98c3B
ge3uWaYZIUEckX3bWgLnPsInsg/2ou48bI+96tGb/agvjLDD1zFhVijQUDwlrIEOYc6gQZ/pjfgF
JtssFsN4zpiIpxFvPZV+ePGc2R0Q8azn3rUCGzEY4rmnxqfNAndMLjIGH8IZ8ANrtYDR6fBriizS
IK0bkpr8CAUr3ij5wZSTHY55XgXHUo4QbV/sL8OeMMEipDmN7+x4EEmkiAmfodQ+8FP464k3CQR6
fQl3J9e9rhduMXmfu08SWsI2g/44V/+r7rQvBW9vUU1eQjSwYMkSFbGxDvDHkXQdr8/f9oRSH41y
ziPHDZ2V06vLDnJIfQ1/FM8OmhbKgoZPMUWAd3xOro1TanjUVs8RKvJSXQMmAd6kC6LXKNmhe7pq
c8YrMxncHVRYyjgrpZhjWCcwZb5e+bTk6PlmgtT7Y6IHtD6++yn0vWgoJhdtW9nDOBXmLENj5mRs
c12lbsy8TZ0+/4S7cnf5CQSjnjKre2pmp77+a42TPEiSGMqnpJTi/MO9NiMzlZeEDgmSVAjm9hx0
HIQ4mS9i5ciZr9s+ibF65wAHO6H72C7wHyQJVQGp5FoMaDHWFN9i13ubj2Vc7KLoWPqi8eYJMdnm
qBP/AgtYXmunowPOvEOmm4weWRluJKu8C2IbN4PchFpS8sxjfxYBMX/g6epyRsRr1DjmlEvUj7ta
WECNhiqx7Rko/psoNKIY1pcJtuJAQi/a5+Nmj1B69tIstVtdT9AjzuI4BmHrdY3TE+qJqMypxRh8
d97hOnBGCChQofLxX/R8x0afa+nOKjp4l7297/byJEqFPtQbZNRCz89eLrIvgyV5UiRvducs3HzR
aUDy88T8+Hax04VTYC+UrqwveUx/zc4lIf/wnY1TCyIdhD8EbTRCKsQybZxYsrwl5wCAnVnx+Gma
fITCs6vsOn1d1qBfxmFY5yJWmzWCd+tvRMz6vr4aWDFl8EKFrx42MUMMIe+AyXzPS9VcSZ+AWgKy
sLVD9fgxQgEdByVymGKc37DJ+81wulbEeUdj01PdkdmXvfsgDrA0fd+IoP6aU3UXN1ve+wnGQESc
1A/qscNU059JiMFUmbOr0GcJnHhsr9T5sstcC3bC3D9XdwAwHx9+nJxQ3Y27CBXgykcjW6WtLS0r
Lfy4YPF8IyGpa3D/JrjUdjm2wTW9tnlnuyzMg6lWqkV0zwX7JP4bHRR1wOXgfbpvG573xe3iUv+L
Kgn2Uv/Rah85uH8bo9EA0YO9IyBeB4avuDJMtn4seLbs+JKRYlqC9MyiqkO/vslgdJ0JriDepTlL
GWbi+EuwrXlu3igGMETOfNaWUM4yDLkWXCdyTYJBTgh8/m4lutvwY4tOwVl90LjAR2jXMCA5csWq
+bQvxPg9bkbKrYsUwPAYoI8q89uDLvaU+/sed6a0KT3Yn0PGXyKTLQQNOh4eefxb9XnjEp34AvNq
ed1WqsabaiXrBJuseyTVNMmSlKCcmEVLY4dn/f2bzMXfNQzcDeR0l3fTdNpre5nsPlEcOOopUvzv
iSpCeW0lmPI4dE3YTBs3ocmEbMWnuohsnnORBtF+XR4bah+WrBonRhCbi/3bFdNEob/DpyMZNpSB
jpUC/g4KEE0ucZDgEnopHg2sI3XzbfwYAI09ijQmBef9Tht8xP2M4ao3p3DZdvK7C9HmNMLJ9eaQ
V7YitBF02HfbkKJHochGCU9BQ+4KKvGovD4dBDGf+37zFgd2VixfpANZql7/6chWi9EZ1WZS6eyr
fMq7vl0AlOCAv6EwJWOqcrLOXMe7/S59B/VzROifDQXh4DiIm/TfVfSUDQrmjV3H++7TAkDwYW+y
064wys+c1UBhhv5qe2Cpvoc0FVbPPSrtsVrnPA+c0kItx+zOywFJMDfO6HrE91RjHn7FkZBMJ2rW
fsy8xVd2jh8ohupjLFP0eUzC6Oco0pNHM/mIgv8A4VYX40+NM6eBEqUcKYehukliujt9DJ/huzAu
oNa9MLN8pXl2lDkD1PJ0//1QE9IBQ2CrPo2fMnn8PW2UMbaswxMhYiTWLfLIGCw0GyjMSibbzd5X
4r/3ZJpxILlTRQUp9MSEvnlqxU9YXqdU2RA4J9KJKuvpMngfkTWMI7O+0HJApJFRx7KkSDi3HvWy
mZkb+SjiwM9TrOzLRxMVkLwEWT+Obosse6HL20C3JHmf50Kqx2/vgs9E1WK5VfbhgVRJLYDyXxfQ
e3gz1SVlntl2j8Xowl+s8feO6vnvBF2S818IIuuVCXAj0jVmzjegpywYyyCWaghK/sdOA0Hz5KPQ
tiA4g860mplfgSwMGK2PiKWJcHJdKkPoZ5ZyqnLpVk0F3mQZG7G1IuKjGgC+iN2AlQ/f/QbLijD/
k0mYlKTXmMzBVBjj1Zyr8frV9SsxOhCLUgTf56n1kbf0YcqqhoWMIoQ7ZtQiBsJL2zVX+Wfxck06
kDb1TLWZDmK9ZmHhq6rfiYnI7h0wyYZ3otxK9+bhkmwEqRR63hLDXv4+uyuVsVcJn8Z/9rN0rWNe
AwEgnLSogNWS/sXjd/+kyDFlLRkniWL5SUCoPXCb0PrjpFrynCMe7qG/cAZQ8JXJEFIEFLgT1L45
AodXf3p0Bq63WdU/AYnWG2pmNHulGrSyJ7xWljJPdvUbKcFGL42DJQUgPUupRlUMCOj4VdEF0c+N
BMh5CF9P+uBSWygUAT6xI8esdWqDfBvStVcc0N+rFwRgscJi3f7lvQadX0Pn83D83OcHD0/Dzv32
PUF351PpVfLT9vpCP4HT3hwZp+XpNVnLes6SfIkgFEXst9Yjtn01wC8rxUBS5vVA8oH3gSRuQ5gp
QEUDHX0EeS+LuaPPUfLVw29RfNjziP1A98CIxq7k0B4HWHzyDzpQp7i0UPdhFWLmOWKMDksXQ+Ls
wuQQL22fv6pPW1835V9FLC1vD68dOjiSDlymZSr32umjb/p6lqB/IiCqwx7rm4q0iPOO/bxkB7Ct
XN9bvRSSmz82d1tuv3jfrp4nyUHpJ7LaBA+JslTCCdJ6Zbz9dxiIoNCYIWi7rY+PPeV7/FGzytH5
dpAsWKIW7qOhEl9xaUDA4Yxy1R5xVmJp4DBgUf24h8fWEOnUSqV/YGvstUv5u+BYLyyP6waiXI/n
BrHCOpWSu1EPG/dzVLuI412WqxnrGysD7J1nQbUGYSJofoz+018RiFRvnp4iN+DoSsmwkFqyLniS
kkgwMZJqjUcX5Bn7zDeDQ+amwjYlfpl12hrHKGJ1SEFjsAElk0azm4WlEuN2cM/hoZNZp4pu2+d/
LK8eIhlOKPewPv8iqP8PrtltoNbf5rjgSXhDZ8Fn/XrOnUJP4CT7KoL8ygk/UpBZPSQLbTRR4X0S
koVT1YCruu9HW2MLrxdrTFeRWCrnq3nhPchDVAA99apIe2A+YtXlFP1f/XO9oaUtFUkhHI7XYmID
PeZmv8TUxrbk0RUYleQl4bW/W+KAZExWpp/ZGZRtgphNRgmRN+Iawqhuq/MUtzuOgStRk7c4kVvA
O4CmOqNkMP01CWy0AOsV76qY5sACsaWQ8bTn2MqTCSVSyE1aqSToe816OolepcgdJcQOb987Gww5
lHraGHgHbo+PaibBTWbQhFiLmxKYdiW+QQ53gU+vQS8z2spEnGOwZuzhI8E9s3IYkfRbVEuHqDfT
YI/XKAqBZc3UgiXnu7RIkVY9XUhNCKNLcMmFvFX3EZM+DchQ31OwyjvpSYiQxhdEK0otIMg/swrV
jhOQqpNgxNak7/iiXwLcpEbqIMxz060yPxOIxSKifVrEo0E4PvY5se7rVPAaTasdmmhkJGlL4J2f
47uRaFcA+SzduZTpKEyH3HlRvx9QvqvIdA5CNZPHX/2S2HUtfsEMR5dlFaUvCAD2TzIJJYlCB84E
s6SiF8Yn2EmgjVByK/ewT9QMK6yWbIQW0Xwo6IKubCrniiQcjoDNKFKF7J4TZJN7QBKYEEvdd9lc
Lt5swBWa/4RgOJ9rxdRBeJyauRG5wEwFg4LZbQTuQR47PH5I/sudU0eMHgjxDhPUSp1iotd6kCL9
eUXyjCRtRlktLPpZeEOL34tUrmdbAtB+YfN6cUJYCmrd3GuyGeup4b2eJQIP1kLOvT50Py6iMAW3
RIAoVwQH+ZJJdTdabMy77dPm0YHSEMjdwKRx5TdmV/gb8X7im78PqOFViSChZugxVHPopEaW/QWz
5+f35HUkwpX+FYOAJiIqy+BHudoXZ+R18un2wosFtciIB16cHc+P/kVDYoZ6DT+7UJrah1/w8DoY
FB8uZqXpMgvOQK9dlr6IXJlwV0NOQOB14lddMwIcysE/rhe+JwWukhzJ3fS0xeTu4Mt4bcCF4KlZ
nO5tyUacAsiNaegc+20CktmLLCKjwfT+CDeuyEHyDKz6TZC6zlypL3Qb5ERoC0Y6dvdxqHA5N4R/
jLN2uq2sL/8lbMsAuOriE7cS0WWYW2ggMqfskzIN/PNhm94m+FUh+26XbcO7jzEkhUeczMDW0Avy
QA96KOaBnuV3PoZuuxlNczvNO9lPqnpLyedCDP5Bt+JrUxmd3ZbGDy8J/LmeGOqTmT82Mtr3bl8B
4fIPzvAwj1W5mrOTqSylVH3nUH542IozIC6qJDxhwK8pngtS/+ZsBFCrPTI5rJIygsvW3IjQVrHA
JsJkS9BTut6PGyWLmemOP7Oiuomutyf7VRKOcHOLXxbBSF78cA2uvBtplDTigXWUvrLyatE0Fw0x
jUJNBQxfBtI+xisin7pIKPjw8v+ghrXp+epTcHAxNBdfjrplIj83S0ndUDarajOPqB5An7tqBU3n
DwYEQ9EnmFTANGuj3XXn4LiVfejLiycuwORHUEfNcahrO2oFou+t0Egi70/pJlCZ5+PK5N7sWRvx
v20Qz+vQ1YziKExKm6IUOLNe74+JmY/ZZvNRBw+TH1ZmEHTwStL6treQvokka0HT2UHCG9ohPjAv
4WfMvvrpUfKz/jJllR8hnMyFygn4sXBxfDox4Mt0uPoowGp383HASsO3isOofB8UPRdpe7pMK5ys
cKEpqwPl+HKJJSDnSU5iy3d/WJBGtUFqHyDFx6qquevprrOijS/SfMJ0cwthmHW03NtJM2FfgHdw
BQ1StCITtze9MAJf4MMof1CgpIpJJSKjuAfDR3l9em5e6S32NqRos3ofFSenclLJylgpqcgsFgea
OdEVWHoS2IeneWUyI9vEGJTxm6B+j2uUCcy0y5hUATYuo2MCITh8o77m+T16XyONVOx3n2uKOTFM
DnHcxmfuJqWrDTohAanZV89WzctWHWWF9Q0HQ+V+taiEALdedXuAFw5UYaAB8/3Yz0pjThD5tRs+
kgmky6pDZI++tSxIz/p9WsC4EkG1Q2R/PxAKxH6DxRzkHsXidiEd6O3PrWj7ippuxqfZhQGjgGmg
CEgbF3Po6Zq7lEXG76WsSZQPAx9HxfI6nvq0I1rd/Ucx889uwuYBFTAxtgB4Q8ajSqVUWS3r9P4t
Tzg/SuphyNksZ9YX0VaVcxOoUsZqIXCCKiaN+mbGUyGi3LwudyXIq9pHKW/k1NE2GiMH5yxJcqdN
YDzngE8xYAy+XV0bocObQ/RWRnKj5oeqMSGsXsXHwBhQ0YeFFIFifeuA2kMC1oXlzIYqVSBHZaUP
22IT3baUaFT0ii8PleP0RD8N1YZ1ti4vISiD6h39ub+vnhGNa22/XIw6PewiSQTGvPu5fRVIAyJO
5M8CZ43d3MN/iDlmnA2VHbrxTZP0xFeu/4OyxPjfJ9sm+5CjSdT0WWfn4usOZams3r8YUzHty7mU
RStJb32hY3m3I/nyvrSCE9S8Xftf79k2TJ36GxbPFul40kOjnqLWRQwp2Bucg6hnUJAJDJnuxzRf
vfF/QzDuwD6GbVaLkyWE27yA7zM9Naj8+NNYCIQm5gWPpUFIWit7rtkAozrOvXOWW9K0/shVmwLn
N56GFxlYS2PAFI9eOYqE4ixjoxt612dVOzR/8CNJosZETnC9O7p3dFBer8GJfT/Kg8Jt7COyHOiO
OMrv7Fhd+DOLPu03Y/lSgEbNO0UUIFymc5FxU9ghNZUnyqEMmE2bH5RnpQUdnRYVs6gitCVvXJZb
/3tkDgP9ACOCYZblevCzaX+9jl3bdju5y+mC3y9Rl9iiyDIQn9gBIeOKEvXaL0B0abdycLcGWsGr
Ntg+hdq14COXju1oS4y9Y81ZJrG+6GJkMF9MI4XHIL+V9bcO6wpQb+l3aLWY0n9ZCnGWDN6ne88F
2kcF0V3JZAwDAbMescRS8MIDb9p5vONrFTAIX7mWJh6R1cFId8l6VXaIm0/Nhk6bncqMAk/REiyf
rMYhVd8zvwkdt0FPMyCT1x5VvjFjnmMZLZZIO666JJkcGXcwN74+HJuUniOE0VQ7cAlYPyNdawlJ
TlSqSmXUi5/RvNAX0cUU4eCnEXUZpySngDAVgJOCVi8sL36K+r6uM/imauYOOJBekXaoAPk9wNMS
KodyVdEhfV1tqQkwKLhTBFXSyB3GMSgDpwB1lOpktJ4QjODsjZi34w5G2FWX96BexaIdy1juE628
1hdiyhOKL98eo4rVqlxl5yUoCXv50mH8Jy1CXUYTxeK36jFhHfTjn9/MixPpUUqJtFmK06b4Fi33
g5zWM4E7I7See1kz4iiKZqWD8rCXYjMqbQvXx2XFTWW/qIqm5sIOtijPISpmkhz2gfMn/0UaU78e
ik7Z6fejBbQ5v59Zemn8DUz3Z2a1/eLxui1hSfCDKotQlkeKHZu6aUTTofcqrEaOjjZ+A6iJqO3f
wFmA8XiO2pGrK08mA9gyw2c9bHj1NPQ/VrFums7eVxSp9cBF0EsedNrDftEuqUW7oSnM1SPoh9uJ
rW8llVNS5q8FyjG2wvYgFJia8+zKZpGhirmIXbQJltYOoy55K63UJpIM4prPCEpAETlsVCbevKKM
l5a1mN04lsu5/MAfYJxm4fjusfanAUWkuPJIj98QbRTgMXgBSfyiNbJ58ONRXLFU3brU6FqnD/ET
Gs00RpnnoCBVsYUJcv706+jPNpK5ndovMBTEEjCVqqJBQcRml5DnS4DtmM8zQIPi3RnkIaT5rYdm
PAyqT73Fcw4Z8n1XJ1xmGYNVmKowuUDOzDkOgGYBxFN0dKfiP+Jy9LzdFL9SIKU/rcKN8CrZo315
MEfNPFIBHUr3cQY9anoCADM6fMBFwpBem8FyKu7mqejJprnttO8VImBlK9D3RKRHCfU6vrcM6anN
LmOxwZXpjEz18FcQysxNVlS3RyHK2u6Rgvpc9WHmj1lrqcOKtIUxwk6zlDriJaI2zoAfZwsj4OnI
uyyK5kctkXSwuq3CUUYtmNJk4xJlHqEW+j0BtmMCPrIUI4D+Nwdm9uo7eRGiVtOr5YyFE6tSiP+o
7zEt5qFyncQjJGtQzblWcDynGA1xb6K2EaE+7uqPp6Mk2qtDGMAZlKidIfdTJCpxNMUAzGfWDjiS
e8HKWMyXiha1MlXRalY6x2tkSJhAsRqpBlk67Wdb4EUqNg1XJiDMR6RqeskJdbc1orMh+bBYU1/R
OoT+oXUPNi1HzfXVKGmDgPjyfH6ncVbV335gjMZJNdHH0FjT+Nf3Xo4zpOipP3eYCnvDB7Gs4vnC
cJChwUtVwdv8ttqk/bsh1OeqdG6NzqvlpKa5aScQEOpKqF15HPNAcvkUvdF5PvcCpERgGUKR42UU
AUm1zKp1hohQgM9Vff45JXhCpfPbCWt4W6mNyVtCmVS1FzWuCuMTpDyFcwgpUyQvsZsQcuAUZFba
7qRXrtBoFJLai6EfJ0cuwfZ0FQbqNACrb8x55in2C0AOfFmUMUnmzHUAMf12x7j/iNT06Jz140XE
nQ6/WW+sd9dTbWikjstNCicpr2ogwdbPXr0Mleyg+SppvoRok9rbd3nrw4DOQIziZhheaip/WNHV
Pu/qGOe/BWEngtTDjNQXx+2gcXZV3CpwqtW3Z2Cq6rY94HROFPOWEHzSPYq9F/ttocOj/CT3yWy2
ztlhF9P0gBrNfFnPxk32M9Fsp0iOZ6nSG+RCIf14kYyFP6YVE1TdpQPRsftZnRdJI2I3CoLCFqls
5t4HJhjhDQm+cxxBTgEwnYJRCJN04U+DmqB/Lh9ojBkOC3zsQwHIh1cG/YyV5bR9LkfXrgReyt/V
OUDCFo47WMjC2unBNfhcN33NUBzp4jcuOnoYkrsh1eBuEYA0iAkBQjmJgGriFINetQ+TQ/z3oZNK
1C9r/T/gfCE9NhIGjNKwB9o0Noy64ZiYUFjjlLOztVLbwPH8HHjWa9R8UxYAaUvEz7oQWxpYNA2O
gM6hQkDYhZFn3PLNm8Q1KbzawHcwQkBpbsccKDkd184WLO1HeusfPdPZkNyp4x4++VyMM+GCQVHT
DZkFc3kA3EJkJPL3wU31Tc//iKNeM53sGLOsUAIAsiLiN04krdFgJ3UGc44YrnqBoz/yOhkQpQOP
km95r7j53et09pnU1iWMtncMQTZ/5u8pEP1kOaKvFlJZt8VRU4hFSKgIrvxTxGt/oMbpA+OXTium
tTvJ3tiLcJOTM5nkndUXeAjSpibiFyfy8CYo6OxAdQiJ+HIHqlIfgyvNyMV3YzIVujGm0j/teOvi
hBWDo+d8IBIy2BFzQfUDYt+qfTm0L+mRo9jqWFgYv3EFRd5MxIqTOPZJShO/rgF0Xt10MP2cIk7I
gp0wiR25ygQOWAmi5IFeb3uabFymxaiqQkncuE6cmkxzon4COniwf9EHUDOD7VNydVa2k9oBHiq4
i4Y0u6k2DahemAqy8fi1m/Xk16HHlsx/LHbPELWSr3RtrP4aG2puczvgd2bLtGdffHmL/QVWiaC8
6/WzXlPSL18EGcsb/OcFBw1Lmnee3O9wcYpsINgX7jbovaS02KryNNJ/ZgGquY0X5xFtoF2UiOtp
aX4giXYKJhVq66gkkuFF/1fvWUpv2ETRFLB9fBhD5eTxiP1u+VjjjeyqeNWIlNMN8i2fRhOkCpBz
63oTf00ZMWpDDKkvsx9jpBp7iEwvV92Zrk58YJVhnRkg1GtGswi1yueB81Rc3TC++cNxOe38Vyuz
gdZLJ3grmNyGI4yELp41zYIWYPBm8HMhY6q7mepSYptA/JsnBZQfl3qd6Bg1WoNu1+ws04UMt1Ih
EFMP+4daRFwpJlb1nqcZZtXy5Yd6lKbZMeDGgKEcsZXaIm0BzVa9/jukF3UKj+QdHoemp84zqFvn
1W5bYH5HjQfKFU2WsuD5lU0xzPcSh+yH5nY8GUKumX9NxXy0VSfOl4COqovnWHSPqZE631u8chPF
qq6+el2Qpy9bLl6wOPgk+ZjpiztgOuCEqRYNbla5jz84LXBHifYc6YNSObEJZtv9VBx0A8dqA0wN
U36UrYfnrNtI1G7OmpWXuaB/BtmRxThzuoe6sCHABODAHzrEY+NfDav6e9sisYLaGNeYnnbbOCBS
FCgu868wti8wMpY4T+vVTzsWoMo5iuHSZz5TgvB9X4qbSwOBeZP/oAKAZXh8xTpyEiCiZjjzL4Xx
2XQ1veVhwxkfcVIOCjLyV1RY/6cZ/E+q1Rk414y3DqIXzGosLqAPe+naa8gDRfudy02EjQZmdfBk
cxrILPqyWlmatwNyitXMibu0YScFVqn5vq0VEpJgIng5pOKrWlMy69ZqciKAia2JqWCdLcwwgd3X
Q7nvnSi+fLTz0gM/FCiIN9ae2cp32pdjmKbmwGUPqaGThVY0ylFrS1FxjUdMLVTbwVK2wyNeno4c
V95P078Cd69+KTMVb9XMYCIViOfGaYIfGixhOUnM252N1qRc8dy35cEoaVBw8VyCYioB/tN/SYNC
XmyZDnj40WMZ6Er/Td9+cw+3W1ESiSm3M8kG4PyRr12GjHBn84lTzFIHPEkvGWDdqWU+q5sl+oQp
sKRI0r8x8625LHBukq9XkJqURYHPJ0A2RM/1nXrZgtnTndDyv8oVQnHm1bZ6mM7TySXU9b9C+L2J
1bbsn1XIpXMazJgZvprN/cFd/6q+rg11lRP29iSc9rRxMhTKggQRau+iWifY//C2JlAnlA+k4pFF
bAFf0DxsnzYQqB2Z2wwsMkoD4fzEQCxujPk0HBW8VRMWXCPtQFLPrclV7InVSkYdp+ZITSeyZ0Z3
NgFXIicC97b6X1QaDbHLUCbWuLPC5JqnCWt5Ud42UMuRw6GITaGSBqsL4U9S7ZO5/6E357X/DWWq
OHZHtNbJRgY0MqVnJ6MowR7q3LAij6q5F3MbxslfLaBvW9IIS5JVhCnKF/isVudshgUGd1F/IME3
RtWXpF56YyKwJOAj+jNGtCUhZ32A/NAplvN/7zsUtrKOTb+SOqO6iCLGgeb5T9zU9G+O3XOcJy7D
MOmXAh+TnzkKjWCw3ik4CCrqPJN6acJGdk2l9EqIdWXEOnHG0yLDFrQBObSF7wpSniJYkrIaef5F
z9HrrATN5FZME4y8oNLj0qa7RTOICI0a9pMpXDbxXCnHVq1Nm0Yjb0/AUv8AcdLTPPtSjvMD8As0
CZJOjcS+XguXERj4q2Iff9eHH3pfiP7Ke43l0HjNbJv7YlU7PSDoboSMXbNibsUAwmsu5QhK73c2
+kZjnusTvI7nHsbvhrp945+CkqM8NWGk67RVX29fQHZ9PzkDlNQZSZYTiLhPI6XxMwFteqcJq3Df
7bfmvUNEprLbG0FAd8xniadL8P+Ae+Wa+35zcWHzwIDrAeZauq92NMpsJjHOAZ5U9kPE1voXY9ed
kq7A9YxUwAfUvkO+CEwKCSdOWDr/rCYK7uqIWzO6yQa6Z8MvbUZ1TL5o/fjSJd0nYguPOlbXt3rc
8yg1VtfI3AwNPfvrZvvPGL8iSSz9Yh4o7QqZTbnVr9lk/FmaiMl8puxCgx+odpIynydkXUitD5Sg
JiShCA1SudJ8cTGM8bk4qvNWq/SrHCk30IvljzRaLtj/+2H0UrP3TBa3qwEN16wsFp+PBtGoKp3h
f2W8xjIBxVqtHvffHCzhW6/4Q6DZrDOBacYwRIX0tLtfhPI4AiZhbrn5YRGl+eKhVcgo43A2DtWG
Vj6ZTU8dCPXWDTaOp0j4EwFsxF9mn3XAzTUnrj+BzjqOouZkecAkBGrZt4FGVqaSuc4NVuZu0fv5
c/S3ugYCwE6kHBK3aAdp9XRNnTwNU6GLKKb37XLZqWWZokq74lg5t3WfDdbqHupm34mvjp0Lq2rL
3TvLB15oGk4msDmukmpM3YQY26Lr67iVffGEIU1CdIvNVyfpuiGHTwk5mw5nDQHHRy2ewYtXW+h4
C9A4prw6NrfwKSTA5YwFd4GiQrTTMgBcD/7WkGpQmMrx4atwSmBN1vzEiN4mnDRuvxSMD10hesTe
+vl24G++6Xk4B3zHvT4yanQHq3YVlVokie35FKmYzYpp6ZYzPxsVmB7HbzxgLB942s8j6Nxzst5I
ekYiK5wRegH8KdGCwkUDrXyR2SHdwb7w4cQE73tRkol67SsAPzBnmMgJq1xSgXlskvTWLeOnsVG0
Y1HU1q6FqHN/ee05QF8ZYWZ7BUVvD8bWOpfk1/yuW3JjuNm3+iM78ehGsLvOY2f0FU3UjlKpx/VX
8WYorTl64aMnBzGfQ0KAQh4nY43D95Ev1XaM1u6QcTMuCtArxsG3BSE4O/NSQbMusPZGbHg2Iyte
zvjRo18cAWWmRQtr1Klp603r9T2YplS4OV8qCOOdGwlZjr4loI8SkBsKf1Kn07WbBv+GC0u5wdlZ
eV1XBSPMTSW8OXq1N9cv69FGMeTiMn7oru27CL7E71zkfOBC2ohE9vRwPBr8toShTCGQVDWFMKsC
3UVYZs7n5oYaKTgc6ZEuqbPUMjKg6Vq0MkIrDoDzWHbJCSqBlBMzn7h/IOEJqmDtYI0WBfEF6GfO
bC9B7DXHks7dGFb388rT8dPnvBHzBt+25Bt3bVn/9VPimT6qpyOq+TJ+vpyzG9V9Wo9YMSjtq8vA
bJszNMGd1a5+8BbKwxjYHb6ua6C5htsCMJ4QTerBn9Zq3dLajZusJif9MNmCQ2zDvUfwPDNbQsj+
3lSY8qSlPGu1fEEjfTXoE2FVX7QGbAnkT5xYbNjutg6psgiwqONHArZJH80fcGN322+Pu19iPO04
hq/HHszzqfYz7Bb4n8rFR1FJdSMYayKPhBru4TcO4qjO3G4n8UNHD6Vz1LhW8nnjKHIklTpPawug
9p2BxApOfSBcGWRkaKSzTzlLQtohCHKF8xyQ5z/cd+jnlDIMr9MQoUSW7pxEKAUOWsSoqkXDysu4
Je/IAJFl/sOG+2UwTxpn0EcJLdC41bYlyoix7QrTQmGBr3WTtYH1IA6dtSCvoSesbPmL3d0JxiFh
AMOHErTnyzc65PuYrM4EcylQZarXhcJZGCMybIE+byQfzWStBqdS5B5uHn36LCRhiZqFKGWucPSN
8HFQY4ksi3n9tmLzR9LE5f7TULg4ZtFy37mIYCRkjEeVwcubK1fTo/LamaikY+LJJPGQoaa241QR
WQMGT4ATb3XNeMtoetGIX7YKJksWROwXou0611q1ejIqH2Q/eYsLX7HG9Z5UtsDfaUZaMBx/afZd
VAzYCvTlhxLnOYJ/KMZ5Z45hyd4w/UeuSnEt7nlkunkvamVMUNSZ9AhO8AA/cUa600JNgnRNL113
o5WqNxZa57HsWLJSs2X17rJplnN2+QV3ChIUBxo9nDToodEwPEKStYMLINYPQzoCRMBOHJa3gCE4
HAhU3LaUXIQMLpgUnQNrmxHgHD5xe2Gj2Wt8DeVCl6dBRFIH/EkMv0rn179mvxrBupGtZ+8xIE5K
lFbbjQjNWH4yj0AlShufnVteWyxSxFZzigNJpdaTh0JUUpKUQZ1ynRh+LxNZMNLH9OZ/IB5Tc7Bs
oStECFhfBD5fQUIsnLAKh9aKAhUoqnocqEMN1djYVALOuhmHixH3gOMQ+KOV0SQASC4jPiXVTx6m
LXZ9ulo3/gk1G0SEpO8JM+nHvtpAsA9GHJsy2HB9cKK98TpiSylWgCSt00oPFlQyQVmvX9HNKxFf
KfRYMkm1KFH0bYpfIvjdBb6ypcBPu+WhP0ndHl4yeav1nfwCo/nHxmsUZUu71ZN8oLdojlJr2tVO
Lg3SOYAJyUzDBhEjZvRi+UexF69svX8bhIQttmPq/LulWGMu5jLBM3gi7gL51iT9QeC0UN4YlL1X
rglmbsGdzWEBAlRDvaAPdY174XiiR+QWUxt60ANSU2hMipNRHvDgoDQs4XE/575Mom+KgJOmh3Le
8fjWymwAThk7Wr85MD3LY8GVuNmrPNNdXgINhwRWakvAT9tDSFoQvVXIQElZQqCrDnaLLbaDJnxl
zfl59/zk6VA63uiaYdtS5RQ5nmWEDCt8bxbfqrYNBIwC9FTEppFyyBIdlmoU77uUBCZS0mrP5oQo
v56cxEj5eeWDD4ofu5P8Adio1btpBRHmwUFI7yJ2AnsI1x1CF/XK1k7lFiBhfu2xV5pYRCpct3co
AkpICuRkU5xxVl6AF/IyrgXnPqn8y8wBn1metDTNcKnTcV8eFsJ2aX+oH1FEcbM42H0m6AYtkIzP
lOno/FJa2/mpKnM5dJNN+pTh3SV1TBc7BZ7g3R0/St3VYEG6wFQ4q9OzJe8iH7OdVNqLiDilouxO
UcEg3RkoSxkS9FZng+K4dfxXCqQ5f/QZFq/rPBsNLZD1iwfGzhGUZRoUxFAACaQUTzZ3qb1YBai0
tA+8zgwDGli0iTlpcGp5KLsEh4G4T0J9jjQ8gJaGlroC8m0xiEJYJwfahSKvRPb3hmsnoQOn4Ipv
aifw+uTUq7vDFTafAKbZ8ju6afpLMJS+bxbwkUxFSjVvnnIZqKMs9JLaAyCNppNw9LnTVSR/4RpU
B90cFMYEABnbrBE0/OqRnM/Bn4NL8NoTt06WIairbMstzO0YtgRz4j/7R1uRNjr4uLVjBfJrrAoT
NTx7mL3Bw4YVx3xwzbmYbX8HkRMuKAVt1BoILB1J6Kf/90yRLitxrF/9kFJ1OwQ3YPEBpKvvcxKJ
jJj0ZxPe6k2Ckaf6AzhL6h+RK8QZFIqBH1XIEGiLYOl1GaJLdE52T58WVGm7aGBeanrM7vLKJ1gA
rx0TfcAQscH3Hme14Ep9TuSSCddmRECZJZv+jC/QMHpoql+x/2G6X/DMRSL6rCIyIJUk42Ktm88A
89s6LhZQdwMgd75MpUSaHbPDoRfS81sdgqPpbI3W+0nUptfWW/BdQ/AA6d9CCPTxQhdUHQrz53rO
EBtdrRpygEId+v3t0nkHMKootjhhRR+qHMnTak5TlPRDWJVxYkMD6VxJT6TsW/1fwoZZsi8SYK4A
PpGjbR9JmrH2+BM0RWi2mUiUypHPa2pSHvaGGPqI4AyJEFM8L5pRRKh0WV+t2dK1WxiQZKUS+qWJ
HMNLsdu3RSUqCedqySVeGP6knAQg74rRXKAbHzBwJJuhx0nP4fwvySIW1PGCpzf4oMDDx3A6unQV
LnzBofeqTY70pHVDi5W/8rFVajfPbNXeoy5Lp97xKgyYEALlgy/t5htGdML5I+iBnRnj62PuRYoS
2jxnd5o+3a0LQW4/NhlZO1HPta+ANrBswmoujtDGCKR6x0caHwxpG35K2htJyIj8o2T7VO1rbBqK
0c+SrEqjexEFoTkiaTObK40WvqpvA3dueok6t6bkKlnQ1SLOyX/08Kv3QqSUNQkMe6muupe0Ue77
mQIjknL7xnwVYyaLH8jbJqh4D9wvaqIbmG77jG1cQauUCnYP5Tt6ueYtJdMaq6xLRNhVIUJfz+d0
RyXWtpfMrS0WOmttvh90YOflN2IKh2s56rr6T5pRZGXSZGtVb81NEsnvJBuqGDZAbq2CubF+EXGt
G1hW/QiTRPB+5RLjMSygNMFqZQbypUlMQ1gJ3Hm4ty0l6crR4MF8xdNES5q77qW5ZgMImNHuisFS
RVMG/4DBEKObF2vHMl+aQSm9SGRQpWSIQzgb39bpz8HMLE+g8AsJZYAvG43q9no+INLvaqfb9FZg
6wkPRJep3jYvdGRRJVFxQQgEBX4OGa/S1iYwTwel8NdsJIUrKskg5xf/snZ0MMWXOgvQ99Wc8yyQ
Ty5gHjbB5ynDCfAyXXecSMYEqYtF+rgYYRmFqwFqtyO94GjwXgw8NnOD6+GgcnRYGLVa5o2rN5+0
AEzT3YCmlfKCw7iFZluZ2yceZcdrgr2oZjrR0fbh6fBb/f40YslBTRfZB171cOhfrBGv85D4uhb3
67r12N5NdRKBwCTIRlnH5cN9I0HFgISDlZgMzKITX4HmM8xGqyyF9DQBQVUwISBDeHx92ESjg83+
mqb5CubTE3yAKtucBPJjuCCyFBIlfcToHklkhFgD3k52vcZXoeQ8JS0LzQrU2gRatLs66oPuJq5i
3mC7wUZJqaPNjNUqzwPZAzoquTp9pAM7AvMWktyLHCtpqH4X7TWMUO17EZX42hH64to6bCtZQbgk
PYeasKcxVVtchbezQMkd6Ok0IVjnlKjOwdbkPLQEBe2Bwwlf6JR0v9hkdWnnPxjziFdbtlQWfr3j
igumxJ3YU5LMlHfcu1Sme8j4l5teLxH8Tjj0FxyrQCOwRk12BG85VtzmBgjf4D1mydO2TcZYUwid
Z9jMtAmDDttUrRa3o7CrYWG+4CZ3G6dlZabHCQlNMQ2N28+sDQVhfBZMEQHPGQT1FGvfMushSruR
4Y/0rhj4InET91A/jeJKeWOl8Ai3tCIIvAYyPRelKBsjwcp1g82+UwZ0pY/MVp2SQJIs9PFrBQNr
Vmy/l9tRc/cya3ACbnL5lS+j6j7eR6rE7e06ZLZqTmNB4pOXYp6a3XADlo7Y4GDP9n2oqS4ptB8Q
p/89ch/DxH2r8Xbn18k53e/9gV1VsN5+hLPtUjPbaBgnXQ/vDo6Lu7dy9GrQId/O4ngrF9vZmOev
2sXxB2799zlpl6WAtPlgxxwfBXR3IfZigYbU5SnF1+IQ4IT914JvF2640iQZWCaDFp0R9alrLzm3
krL/LlInw1387ZXqCM4u6DWzv/zyEEYvmy9erodvFxkg5IxmQWziOwLgR0DQ1IdXzreWZ7adzPty
yNSi7NdNK5zBeQiBMoQDrt6JK03XWKS32nMtxcSsiEjaJaJmlCWdCZDwVt37L0MEmsqR1nWfLsv1
qDttyNHM/NDntcc6ybwiVhfmqIind+0b1qixnaWh52pecGpbUroeKiQxBAf75Wjc0ZOE7f0/D7J7
JRovWk2D+fpxm4Vs+FbvHkCKEg8ZUhJGWayhUNPtjHTMM8Z6mm6jzPtLwqZp8gYr40tMjbi85MCn
bg7X8Z2nMx2i0fdwhM4iYnAFY6J5ARlWfgP/jYmJDQpMFe6DAXXh16n3O/lshV9EQ/vbG810xjD6
UK12cQdTx09KDrXt2SvAzzocPzejW13H6zSX4HhkjzbaXXjVrXQvmIvq7+b22q2L0Sjmo0AfmsdL
OJ602Ks2BY6OQdlombt1NHI5qY76JosB2IQXfuwkHPdY2Rw4PkVznnXQ2hrtKaHpYS435cn9vKbL
y36PZjIM/Baa8kbn1BXsFchllmsed5C6Xq0oSSNmrVwID1L0Z0OsBhO++sjkjEkSNRqKxBJtefPz
2bvLVoZRdeCLRvHJrpjyqKV24y1wRoaODwqWbg01VNdbwT+wzHVgKxu9sttzVBXTj0TmdebvqHns
AKyCIsf15dADHwWm8rBKFFxEPii0HtyTTbre25zVrsTCtsKARfcE9dqU8hvd/71ssdLfbxVbVCpp
sOG7B86ffC3zKjz9iJ/IbEyMASK6wlC6DNEx2IWsaOHVPo8Kexcg1+miWAp5pLM4kxliIxE/sJpz
fw91Fh4tNfNTfCdiXGdZJqPAl+A0I+rQSyHGsYZ2R/lh1aebFD9t7X/oFgp8kO1iScdJS9cUwHzj
w0TLeXAkfR/QijMGWuqgKDR6tDj7HmjMv39rYCFf1Bo4barGURAp+KIAPQS1kx1OpaZnIwJte82v
SCiYVtJYinRwqxr2eHV8V1PwQtehaj8q4ZDllctal91sCexXauwljX5bNzr0U6qNjRDwf+iXvCE3
WvsVuCY2TSSGgc6pazX7a+Q/Fkzxt29tVBhdXLAjNTNTEfNNmU1mWQjLYMoWNzNjxmb7qMYoL9IA
uDp2cYvpiYed09vkecEnYOgMC21A855UI2PrfK832upCwqvvCQ1LDoITBJFwfuysoe5hnpmhb8us
b+z2ZOgTm7i8AnQ/Myth28Oye+Hm8azpU7RxVGk0pMt4EYnVa1bIhVB7ClXV7SGtiD6Wrkg966V/
GG0IrK/PGlghucAwdiSSzPbKbA5ryX06D+W/FD67VWGbKtGouq/I8z+CSBys+2hGzzNXRXW91uKg
KcLSKKS3vuak6FJBz/EfLQaDd9YNcF7ZKVIJCIK3T5QoT2B58xZmhIwmIFGeBK98SyOy/pQGKNCA
oRMKizq9LvlzBZId58+BYd+EWMlsR9y7Om+QutiM2rbQyxPD3b6ddCzdFy9Q07dT5Naw/aNpWNcc
D75GmCDM/BS/WcE9Z4lFQs7sVTBYfpz+ehw41h25UJmxGKpseJVMyrwXakIkrcQAEEvetC9B2XWw
ByjCWL2hzdJ7cbLimMkduiUxfrHeChn6jWd4Sjz28ofjF5hn+jCUI34SfUAijtgM6oxGW3xMI9cj
iK4STQi3lquajBlZ44osQGA+1HPvRIuN6I34u6WrhJwxLJakrbnhH/axFBs2HByeV7w6H0AMyj26
07rSTZ3HYMObHNbfpdp1InKxgsZCgVhjKu94VOOnd8H9t3Zyh0iaUPL1SwuNv5BOBVOx9UjhPCzY
49OYmPucDpTdS0xAKjM4y78LNXmdICSrpY7Xup6MFYBVCFSWu/8bK534xoupeYbnefbifU1XD6hF
tHvNLCXdpFmoos1jQUktGbw/03ISpZvywwaP82FCIJGnvpLpTqLTr0aJT50UPcg0u+i0DVhnrb76
9GDgNHxPrc+pgerHFHH6JKJfZpVdQMvaIZ66lTZvmG3ID0ctusj7QjY3g9tK2gIJF0ZQuu75ems1
t1Tu7FREBKdDbVJ/TdxAxictAo4fVfeHt9cbmf42/RcPRymxQ6bVqWTUoZX1LnXjUkTC6MKHuYyJ
OGZWaFslBJ6f8NQ6Ghy1+6ODn8xqNMYRsrjFw0dbCb+205PqG22Mn84GmdQ0Uoqf5KqJBmoSHtGW
aCVB3YJ9v/DXeGIxk+IGdk+BDVhYic2Vuoo1qkHpwZfLPl1OJGSJbZZ8SDE/0AEiGtdif930BW9L
/RjOhLV92/0c+bGHoWj+R8IjuQXvgAiF0cV2qSkekHpqMjK+RagfyKjTCo1oFdOSGiJoL5tzUsk/
Ss0ThCDTM+Rg+Tj4PlUp5LH5YmDq5B6uB4VmWoPzA5O5sZ6fH4gEzPlU0uCD7coNmdyCYKP1cjuq
m66Vxa3CQgMXlmQur7dv2lBaQwgAg/95HohQ3EOVdoN6aHVvuNz9tn1fFnaeKJdNaX7zJ8EB8Wxz
Gebtzb/GqVbWHso/vvVUckyCqkMyr9EopV+QlND76eGVYr7hQmUsyoK/JzXrk2DNMQViM2KmZuUK
Kc7Lrgreg34hBVeUHMZ10lo9RA51Wa2b54ty0Wjcb6OdcSSeamdYS6XYbkGcATcGSMY8HIH/h0JP
Dan6469NU1Cu7Nkb1aqsUyx1HrzZUGkTIutmI+0MuI1wDGbdPZSBVDTZYoV6SHMNXCuRq5ayi72W
cfR/+pRCt3ZpXMAE9Jj3jJiAzVyPSA6SG4/u7l+NlMicafo+jpwoFTaMUOebfNimf3aZv6q+44Wg
0FW3LNOfAfcRXjafl5+F4XPIFpqDBWsPBXcOVE1jfkEmTT6+1bvmK83/5CrkmUMAjeHEITHw8CUl
YrTgk4pjybZC7NpiBVJSpO0mI4cYn8h/oZhgtUD3E1R+rTUDXsi2WqTG4ULZseThuTayKTbei2pY
3OMByzUV2JjVRRWRK6Waff8+/hlZOuhFPhrIQBkG34W7NXT65t3cfX2A5E/f6S+QVIV05msUNnMs
Ez5j1+t2Bm632bd/UMGo8wBv6bRh5JzFar5jBxDxLZ9IXs72wHYSE5vQhj3t3DUXCultGjTngvfT
l5/TD6wdRG0/t6Rsg7XWn/aqslosfU5BVq07iCITv3Z/a0Y8VAXsU7eFQreQrF+0+GCTFnkQtQlO
/p1zjr43C+VTNt966vtzg6FOfamrO0YBbD3O8pVDeXGJUZLNXZtZ6AxknbAwLDPj07IUSyI217kh
oq6bACo64FCIZ+FN94SqdAqpbjEq9/oPm3TI8pXIuNof4elRFoln2+QPOrPKXZh9pCMs0OvKLyqT
rAp6S1eTOAtzL/85trspJy5sr9Yzn1CTSjQS7uqet13VLoR7KuKTQDRAWUHOdv2whyyyEj3jXXy5
eIQyYbbwNQtAqkHzK5Iu//V6Cz5QbMjXbTc18Gijp/xHU5Mk2y7jAIFx1ZLrIOnux/RqQIFtfB4j
tnwn3xJBu3PuxElwbKCxEKgoEDPCS3T7IIEq9Evi7bVAIdReT5HcvW1i5pjwknb7jclRJi4DaM4p
sA+8TYmcPQZt2iC+B03MClg3GuPErfw+6bb76Dj64labK5ydaYbWIddusWbzxVXURFcYF+51QEr9
Z2yt7wNvhPy1dOWrHm4ontg8oGvQgmYKPqk3IbdzC45tNdIk7Iq60l9ogxuCkwdxm2+ljQOpc2wI
UYeda9u1BJvfrTDwbUEjj2ZnPtxzzEFgb5isIC/vjq/xjzkaw1940eUGRuOhpYaH2UGy6GHGUwg4
29+fGt3iXD+12XgzVicsIEeyQ2D5BtcqaiQboD6vRgdBmEe1on2j0U71m7ze1qNqSAFNrI/TNc8r
hZxe/chLSnRsYjktXdhsNbjfL5FzKnzUq1tbcBEFOEf79wuo3VOIBLo2Q/VJdhQWq+rV+pLNFnoB
faqh4bOKCPclGqhnKS0wgqc4g7f5aDKECygtthn06B4LhLXad2chRIeMANrOngVkvfIvtJZq40Zb
9+vtr/uBcUMQXsXwX89eKY0xaFaAgBmmDilE9UqKs20P/mlPdpb+Tha8FY/lcrFVZjgFH8YumSbC
qrNlGtAEZjyRaZlVskIyPiRjKwkEiuZbXd7XGtarKSvdlVzlVboinNcWATVR84EeTTJJubnLUI7q
VjpMvCLY80Nkqwv5do5dSL5N+DL5QUG8PQ0YEBh4fsuaPFB+aXxgR5bKNj2hGjoPbSRFZthGyPcx
Wy0mX4Tj1CgAjVlJ+97czgUUFuaQ0QvAsyAwLUuWwEFXR3kN4dVv8IUdTBe39eNltRW8xneRMuEy
GsK3ahX6pTYHBDxNvp0EDNxyZLM8rxIE0IOlfYGbHUPv+vsR9RfmYjjAEaNaN6evlDTxeRX6r4a1
82lsjhbQ/pAlYvHV1yVWxklORZJYyx9XkwTso9PHuUVjmQNDJ2dMLkYi+OY5Oj0UU1NxSyCKPoZP
rlS6xRQv9zpnfgfWYjmMhq6fG1t+SDjlt+r8UYy4+k3aV2iTmqH1LwYPyU3zdyAJNBrBOWDl/vxX
z25i1KR44eDuN1FI7773DOA1EeBNnA5kS4C06r8rrHCmy0Q4fDMVIul3G2PYZad3Lq4QrKBOoPyR
/vbHW8jDR+tEAYe2WoF5JLkP4Iy8/5mM2MIn/dBEhLVtcnGXMEYrRFctDs2Ub6gPnJ0Kx0c4AHgF
R6uiGgZkzFv0vN5v3mOXLj+BBzcJVKnqTQQ/1vu7mDgzoN4rLjQw5wJcl94nrQRmg6E1SG1uwB0O
SxiinHQRTeaQZo3WZY4aiFool8JS0KkebaIS0gK0q47hSAIZTutf6yz2WXGKk8YeEFgMEISSdnqL
HmNNemcgjJwHw2NJc8JWhqpCjeQqbHQEF2Yb4MD7pnsCCfZolwFjanZHC5ub3ap3ZfhJZuRiFuKE
6AyZp73DamTzC+MAEjz3Rs7Kwb57q7Yc9wxyeIq4oati6zdvb2jR+872f2LplDcQnlRcJV0sm9UO
vX4C+5HROLyDyl1bENnHTWE9oLfg7b0RAz5kyvJOjOfxOy+qz0nLkvIYcdEMSy/JS3QJt+J6pqQb
HGo92OPqvMg4a9w6q/4d2ywJl2taqHp4fK57sF9dMsww6UCfGMc135zpOkPoQ3jDYZ0SbvNn9Cyr
0DfNP03nkcfi00WkzSIL+OeDHe7Ah3m3Juks/JLs6yzHDojDtztozXyANi9Hp1xlE8TgSrufWDMH
tTRN6J5vNwLimN8Nz7pwExR8rNR7FzTtmSgIuFbOHIMn/hAsufoS9zlpd/Mr/MjcI62la19CtrNj
8XUWTMjQ8C00mZ1uIikpZ1MDFQHs0jH7cYdPwMlfZXwToTW26JxFuQH1zIqfItDpuv5D91xPJsW2
fH8dnqWsMNye6akNgJVu2tiFZC18UXkOOkPkpvBxRtTa7iblkWfTPXQewyr4KvICIA30OpXE1Ix6
8LvgTuBxWzNjgZwzf3+TtRX5KDw6gkcGLsLmAaSug2KVr6lBfoblO0wKQNxaY4qGkPjXzOTCgdl+
gSJlQa81fC2gOIFtqO34abcX0DUyuKYfi/qagtRRC+P1Oe+yWXzwFYzkTlGOin8B5VxXqwjeCi42
n/kavLD7dyI1w0AAA6wUiZPMI7X7+rPoCwjlc8jl4AgSW1gePBNRMi2Qso82+LbraoLNdBGf2I1I
eSeQFeNxZHR313mK2xLWSRrv5ErgzdHSKYbeB9REQiN5DE/RtDzZm5xHw/xtKnGOeieEhhhtovYD
lBK7enf+B5EAIBLT9hrjOylb0n8KVWhNeGB4bqSV601F3BB+Br47zd56DuEIfknfRzZ1CLhWOrEH
vZnKAGvT1gGgcamDEAnOeX3Moo5nkdMthUrJaOVxpl0MKh1lA0tSBOCTo/DDaxMLjTdPlpxuXFr8
fszpnu/9iKm6HAOLBDZLW+4je0SeLU8Ne5OgbtwUba3dGl9NR5jsts9PpTgKmOzj8higroxTdQWI
wJlBKAypqrjnlRmpqxrhqy+knfaUuc8cXcfhHPWWAOQzKv0cNXA1W7O226pInBcKF/X762uooAql
EIjSA4LCHq8hPu5HCSx1TywbSo01N9eO6Ee1vlocDOYm4w2PaAlhIpwnBYRjCq8nmWVBO0RjQ6X/
M2WmHf2fym1JOtYl+Qn06Wv3vkAGDaWG1GgshJXIKVqRkX1PXqcLJ7e9P4VNR9f97fxsAvQguSjZ
pw7/U19cXgC99W3RnRQr4Xt+dwweXe3YO3oir0dMMml8m5ceMOoHT5a1574Tft823mCWu45RnTmw
nUtGVfuWsqRXK/uK2yzxGAK4zE9NqcPueYgvqH+S0W22N/Z5AJkI0odsv7e/JMfevVIwAeFJ45LU
brb/C7XKmj9tVALVVDqL0neBxF4zZJU9hzcZ58jQkK8ITy0F1+gQSaBOVZd8y0VQqBghlQNoIguV
eyZuaIAu9AVNoXqw6VLXtIOP9SjFnH6FjVWgG0WRjIRAKsqsh4nXrHDim3/XO2xZN3QuSFDY+fib
NJV44mne3pLCPn+kkXk1CQqWubkWutQgKExT2DgrGm4lZ6kSsYsTAuyajaS5ZVZvzqU/4BYIP1bu
RMay5V874OaoVyyR+PSraCpQbU6ByTPK4DGM3aehEns1dl2tu2Zjt82pCgfIlUYWpHs1bfKyGj8H
ufNoaVrCi3TgerWn8ORSTijwohWLk9xlVyqqdWghcvEGdACI1/9OcJseg+OL/j+YWZwfJMHei/1x
nSkqQkX79QryFG2gdGUCMnu70iFpMbHkAuJpNI+74UJxQ0zj4dk0H49oo/5bI4anGU2jvX0tiZ8M
sUO/m0V6mnhH6njB+pNw0buost04Y8mOsA53gOJ6woS+YDXiSsUtahlmZbxvn6sW0x/fLe1PeVzu
JucC90ZQReEXHK1pVXYcud0U4plFbEZo+kp6G7u50/WppEGQsfy2d0dCLfac60GgbhHuLr/4xuyS
TosMQHQW9AoPp5tE04GHqiY7Z1QSG2CR2A11sYC4bsF2jTz4NSy/iGELsjCDbetc13sR6aOTAl8o
q57t5CWg6mSexCvj0ELrUBwRVoiJSB8/vrULvJ4LOAUzI2ws0seQpmNhPKSSUtwjC8yVCiakuXOO
cirnYUSlNOcczU4GI/jDl26wEVXtVtQO8quyQqMI5ljt4kfxWzRxPupNo+4pOtHuA0yT21m0uhnK
+Pe+b/h4NHsK14/sfEKBGDvcOisozqsAx2hyEXbnHHHob+mdo1OpMN+0e0aapeXtXXeSNmV5U/ed
fQM7hPDjEWok/2jRu0EAa3zwNAY9hJjtcXY/ytLro8TC/0mJMjgpGFa3g9QJgplbzCyrZnjpismb
sqbUDq0nSEvOY9qezIshLPdo7nzeFTdKkIpTZ0uZugv9BeEEnqB1oq4ECuSSMg7bqcLZ0D5iLnzW
yPTwTucq2S/92Ecbi6A3RCWgLKUq/kPS0sDQg8xLLm3sCWtbeYCPaY73mFUqyri2cPoosIji7fsE
OYD5hQf92CIax6wokjafy77v9lFMgr23SnUngB5mcR8B1l5kJ9fGu/f6++o1Cym3CWprn7ntV7Of
RqMXRfisAma3uh+bg93n7ZJbznYnKQemLElC72XSj0u5+mNU1PYP4FuorbRrtIMkyAYy3ChpTdB+
Gz+sVm6hsr4u3gKUJzwGQQul710nhlcqzp1OMzlm65o/nSTKbE7uya73S1n/zsxgHGFVL+syJoMF
cp1aepCRLIwtuovUAsqlhHiuQ9zGSfnamD4jPEfJxCistO7M5jNNqDvXxuvtUtnNDqks5pC40DJD
q5gOXHHprpT2YG7x5UqF4kQ0YExUAnZHm6dXojjIcxABZNPFsjdq31azKaQ8IGnhsMwm9/y7/GT6
/0fLMcz2HDzRX/ogQwwBxnLqnUZdNOGE/+Olj0YbjLeLGVijgR1FvKDKT5e7kmIn8LbwACxDckK6
uEcw0Vo664VKc1ra9hHJwGkjNa29aj6gYnt5CYYQw1gF2Fb8/y7bZJ3kWaOJQp9l3URh5xlbS1D/
Wu29HwrF4xjmWpxYmkriBVh/i2dGPx8qYBcNE1mKtl8+k36ouaUK67r9KBzRCTrSA3EQvRLB5h0o
d5vKyxK7kknWUTER5kjv48cjPI3T9VSuzX4DGp+AzhjNGm+LNxJPKH4ixt2wIZBEbl//69D758ux
N15rEGJLrAnDfA5iqnS4hzCUufIHYDX9quRdbQq08ThSFcwyRWE23lLbM5tz0IbnL31306alX3m5
tF9a3qex1AMdLnBqMOTiMysZPJDYr92pZ9QCd0oXDkRLvAh2txTcEpFT0pFeuuUNAdhjOLe39GLj
R7bIS7AZWJUglGpPyCgzsN7pW9z8TRauZD1VVyC8YdfXOtDyng5mLZkH/MujuRhnfXiP3qO1XOnY
lwdeXSVMEtMFlFb9jKETnQl+VPv/39V6V7StGd60kEjXGZWeQ3FOFVMsRwpiT+oaWyTmEk3i9iMZ
3LR/4qfH+JfjUJWipVGM7UnBF8CYOkbCkb1Mtvvtt40j4sGOsLSZwnpoJUPZLCXfGqIX+wB2ghWM
Kg7nMkM9dPeP6f2lOf187g/KL0UVzcBwYz86SKzynjoaZSAKcASBLHU9pSS6mdN5EMMNCPzDxAb2
dBkiohqQw/QxmBYxkUSSq8/NCVIMQV+wHU4Pz04GMvtteYFAEIOCExtmCQjQ/UFL0sxKCUP2dVXp
pXIhz3WdSU1OYDo2tvj13x3k6Vdo8e3+EF6LxY12Vf/+IEjLFaltLU7wx1ax78LkoWDrZmHNGq6F
F1leVv7tI6shqMHepReAlBDc0Flk8snJa75Fr3fbkfl1lReIDUnTVRgveykw0qtteuKmxAmQsLjr
BD+2Q1Z3L/J+sfd/6kIPcgkLab8EO6lmtJjklmCXDIEiBSpqD7ynfY1JPn10piHoYVoouCsEYCdN
/Tf891Nmvvy9cXDLzDeUCTre3iyNAIGSbkFqbY1WXPpaqjEnHGENN+4GGk0jvszmGGINaxv/x21L
IqJ7zxjRpqznK9BDZKhFuCuEn81Gge/LvF80CP5jZP2SE4f6b5HywMoyE+RPaAscsDm0eAt9g4BR
3/Ca7+CkAshGpdOiC046gkuI9PpXiKNpSE/XrwIjbnG/0y8WypR/EJWo4tYOzMceW88amm1caXvC
VBG7rZ9QhhTOEd2LaFs9hUxAzDQvKXNT700tfOuiifohsfLTOrbsyjTgM6ifHVY9A64pBjYtI+So
0mSaQBUQvsBeTqutZJVSbzr2JUiySHKV+DR1bmn8sCfCYNkdhVdUyxsFr8Ay0mnATLYtfG/CDXAP
ZbZIJhcyncmsweMa6Jt/eeRTMUs3E0Kz09PzAT6BXRegXxS/v7cRi5WsrjdtnAoARkNfNwAZ6j6p
JfgkQYDG1JUAX16o9kh8iVggXazlW+WXI6EKMWJPVilNNtLIaIyGRfpPo0WMFjj7AytPl/ICTzCF
QrwBLpGqee3HKelLkfZHrnLW7+05wkCIhGAzmZvmEUzodxYtNXgaVvEWCshZne1uUyEUylt8cFdZ
uNd0S4Wu+Aiq517kuzCmjsYhEmoupAPxUq1NR/6TVm0ARv7xDF1Q8dpiiEqr8FeHrD3ninMrVBZz
vbFT1Ec14WsefTPIE9DUYn9T2l1jcMH6izJ9UA2DGXpQf8be8z073fID5ZhJQhqZqP+rE3/uAaof
sws5/IfA65vfIA5iVGcCnBh8TY5JBAhjV1R4MreXM5aR4sOzz06VffuEyONRcY+FXPxxkwmjcMkr
Blt/lIEgDkJvhq3lVpq8kU57kVzajvv0/Q3rM90EUhSu2uFWINOvLo8E8dyMmLwkdRtcZlSjCc5W
K8eKki1Z2CTPil7QSY484lZVtA8BAWtPEckr0FaRJdFSoVmm39iBXhzNDjkNLYox1iCGyoFDCFkg
1ApLsT+TOsdvOWoW8+a0hzIDew5ZBWCs2yWRdDNAGtrFm9KvU7Y9ZAVCKtaUKDblGyy0xXLh1Tps
DtTXDNJrmm1mKgQBEBRqmqXE72BkbEaCmo80SFrEwXMwgFb3g1eCVdDD35KBCGgN+56XysTA1lM+
j+UE9aGO5PjYNBxGCTljdNALsqjjL5HFc1DTNcN5SiiqDuyT7Jljf90p7qEPEIWu2rdorbwwY4Yn
PwP797qvCr1eu0Nt3xqDKemswA+7t9OcRrkSfG7q4Gs+1yhevrbTBhH5uHufZhHloKcJWrk71s7t
lqRVAArvcktD4kMpaBSg6kanZPN8xbGLqt7QTHTFEH/4AgY3Ysx+Bo3//TAfrvLvdiQ53cXmJUAB
AWzRJTXuCNVB3/YavyItuAtUa2kl8zPLPEgZMmwd6D+UkR2sTexgAloGeVJr7fIjzO0dtqZgNRTt
J8/iXdwVT+NgbEU9Rfj0CHekXI5F8eUYoCJLYCwDhgcU3i88mxEdoUsWrN8HeYbVG20AUuOaj4/S
GwPhNsrhgLB6nqCMS6bYuyTxjA0B0yRMkuTaVm5EMY2bEJWhU0V3auhpcohXGlH00U3SP1DQIsP+
ENTSseBPsxYahBWHdeXkHXqsbsgj38/hLjdk+WBXHU6Z6UubnDWKmASZg85QifH0THgnn8ISm/n2
gb80tD+92A1jwNrh/rrMjYI7U9RRtS58Nzz1aS3FiqS+C1j8wisoHDhE127+lzfvJQtiBm+JeAPp
Gae3MkFqyojcGa6UPsQBrr0f5q+g8D2X1ClWJN699c/zHZvhMBgNwAHWwS25lbvqs274i/05Em/r
tbNu5OCoC5OmZdn2Y/zbOs5Xugm+DskY0c4me8dlmEf+qE2CfZcHCfjIT36hFXXAxnGq32GzVjq3
HntBh0FUBGH7ohSQsKO2PY8CViXT1AdO7O4zHENT2UZOPntAPVWzs3BR+ckr+zc63hA+s4ipQUbe
jsn94kxQhVSJaIgHtxn5wkcYARPg4JF1/tZzX+8vtu6KAmGI/RCgQAC6k86aBYXC6PIInD+7IKEP
2mTtM5+VS9zb6V+t83KPxQdtizF5QEKbZrMUxgI4qf2m6OCvoL8efcbNH4rhwDnR3ViViHlzgxj1
b+nV/Vk5U0taXo3euZh6ZHiFIYqabHHlV3pslL5VbuED2w40o5dHYRNm1ywZKij+otu83FFkTVBl
HL6lsMe6cmyvScA3JevXQlYGn7egltJALz59VCyqUZkSo7O3UHaR3dUJIlEeTijUVDSfXJSaSULy
3M5pSQXGvCFhOe9745kv9xF43gSphy3cw0bmCfj+LG108X0FqIJ/vc7IdSpTVBqFwfFZbITZrX/9
HqR2FQZIPGKHKbZJQ+/SSVog99c1Vl8Rt+vaGkCyBu05j+gg8lkb+ah4HTHsHnhZXrJbJwJVW4yq
elZ00BMvRZn5kAPg3k7cDNCVzQ3NTRy46UtntTwSNzGoQcdgh+0s+BGtM9VqhExisw46Jz4VG59e
sclsK49qkFSOFOV595d2hUvwYaIlvetdCK4kOzRBD7sfdTa5mX6mGPwdO5M5x0FPUYh226ElxU0z
PjtBMYFWjU8WJXhlBsn6DqOUOim51QLPp33o3Fu8/K45/ckbuSlnVstMQyT9ujKEJ9TPY1+ZaBCo
DtsUvEwcabrJuUcjnCG9MvcROiM0NCCYFoN/iq77Hflxwa41ZnwCrv/6DSEPC53rJ9DJc3K7D7ht
to0k/hcC/yr8g1jBXrF6fBJtbSlWfKILttxq2gk1pFU8r5igoVPULq5vshFhS04/rXKcuwR3mt5T
dGWNjCk9gZmLfN3t6WZWzXPexJFslnKcp/FtITRnazu5k1lubERsjW9LwnbPb4/AjQNmUFWDA+F8
t27fejzE6MuUidFwRlJLFlVRMcjPUB1qPmuxwxUok5S1ciDRHYn5Lw/pc7Wz7cDEwAm4rYKMo3X5
cWT/2oXrVvp/bha9NM82Lbw54SDpUbQslGoqjjhQf3bmZwT7wL/Ofjo4MMhqE3XYkFvEMhskuPRy
IwFPHKGttxW7oKU1a+u1EMvXL8jCCFkNRs3UzJLJMOUTKG9rnFHqCG52oHqh+AN47abGK8aydwKf
9TCEJgSg6KFUX/p2dN2BvUei/bT1Nq48cbFSjauqcoE+RL0BS+0HZKyevZ9M64fFs3/fKU7p3WFd
LLG3rE7BC5Xz95/29Hl+GnI765eJqeyV6m+1Lq4VYMMh6F2agBXxxjri9KCH3KQX1/qhLPiD5uJg
m8emehLZldZMin3M3Z9bWK+zKv23WnxwdhZGvdHo9Ny9W+egzuublfqMqXxXaip0xCGeGHqpgMWY
uQpIbJKsysLgdSCB9wjydjlTHEoKJbeSjGmD3VueIbF5hyI7lHuHFHPkxsC9cHwyLwsjrgJMXgmF
N2kXV6uS7pC44PCezGWhppTGwvUfJ83Oj+17amXxT1vd5CabxedOc0T5dZFC3BUgJrm6JSZ2xtRS
+ud51+3+zbzK3vxu82My/k7ic3m8pRSEcLGoA+vwyB+OjKBPxTu0ZAqGN2vIPG8c4Va7unYWAjf/
FXogKKvcOwXksvftx2pj+ODWAGQwCYzF1FC+Rh/XnD8j8pGefOGbExVKJDVjgGE5WrpiYeD+LrEo
DdOnS+gjCfy6cmlstJGqV4JveeN4xDh9Tg7kKEeDeQclz8ySwdnoOUKZLx/oE7PcIL8ykk0S88OG
HSbhitHquPzilFmNNmeHZg60QJpJ6xGJYRwzHhaDRvem1o3hCbMxvbMlpe0YFttJZkrMZVyJSKXv
A0X6jLE9TzHNMJh2IYH26JujRlz/OvT3B91LaRepHWvJ4MTeSisF6nhzAMSP836/ZWGFwbREys5B
/2qGFsuMoFzTaBKuTAOtj7wUOSITDt1meTHNfYZvy+2fUaONryd9x0e4iZ0E3U7xxhTvUQAPqyUE
jfi3JSIi39cMbev+EzRlwrlbRg5HY9Siom7qKJc6vqY+ErFB6a4EFiXxo8ByQtrSjeDH2IAjp0Gr
ONdkF483+rND6GW12qcPsGac59U7Xu6NvPdaR12fvV9+e1q/kmUmb+uVX8L4MRR7pMz3v+Fq2EdJ
Zfa4nB5XZsHQuJgr5aBvywK5lI3o86ek1ymMMvZ0jJ7x5w0h9ntbqIsBSCR82mnaMviPD3zdtJtr
nQWNRvkny7KhqlopiIZZzKaUaoyBNpI/hF+FAryaKcWPt58LjW/BjZEpU7FG+a1RxTWgpPdgtLSO
AzCsxIqJhLR6ePDmGF36Z5i/BXup3oVZeTNm3ZzwL4mO6Zn1GrF7CZFZgqlVo7Ugb+ATP4fXaiiH
qBd6Z7KZBSs4N++NBWv0RJEiWUI9hIq1Kfa2pEAn9RVwkrwkJdVSZJryC+nV1zUaVwVF5VAcwRHH
E0l8QYxEeXgpo1N3MhIECi4TCljUkI72LZi4sWp4GQOfROmhRCw9HxVpJOizMkh3hgp64mOVchHP
UFioUnKY9xQPsSGKTdlrPsxkdFcMeKg3rwiORtjJdtdZ1QeutnRge6CEG8Jmi43Tp1JhwTwWMIYh
AtJ1mujd98WFj7TDmirZYJo8ib+SL8ss0rryBgF/BOWYfTlpxWMP75LI3AJhxCrNaPSirDZnLNh/
8PomZM5U13VuQNQoxIfILddw2m7XC1SFGYMRBox8g7+6OzX+flzt0NCYJQzuZGkXZC7E1rCoyxVi
u6Unid2MQ62x3cW4pAt+wLQuOOAi4KVD9BW5xKPwSxbgm67Z9n9Tj93IfrHylqAhVrTRksKirSvC
tjg8+Lo3xjq89TzEmlhkFkbyY527D0fqfEkCFtRNzzespLEpxmCMaB0eR7tCAVCveaKjuqmcZ1bN
S3yIZ4nt+DB7nsF6kcShExZgGvNDX0FLnmaXSOHUZujn9/FxFGqCsfzgLAZUaxxbLaVeJHHqHAVj
JCQBuHhVkv5jJj/8k6h8VrCyTyknIYdOGuYv9iMisIPZ/FcPYRmzMVY1qxMUzuHO9OEfCQfEfVET
DCMKpde607vhhxzIAX0sHiphEn6VdIA1qUD6N+7Qy9VEfC8rOQ9N6dyQ/SMT13H3BQzV0kAnrC3N
ZW8rHx4Q2fHGEqB8a2UWKuWzAeHhTE7736MIi4zqhxPAZ2nq46JGWpeeII7xgFRAyWTw/q8ClZ06
UbeQKjOMZUI4XJDDS1Q84/H4Gpxtwui1gBnbrvw4n3j+FrozkyJiS+rMhsGZBtlCfFRYaqD12vO/
u0oJ1SOrP4eYQIBFiDc8umJ6fibPoZVWVYcod+m5MDbwslmHhbwBK7DomECSBpfGHrSUuaoqhp7p
LeBBsOFjqvQlZJ71XqOQQ1NXvuahI7HQ0SjFSMXaV9/6wtqvvKJCzqXuGGrgtXV2xl9Hkuxi6Pty
6t+nJJpXpx++32zsL20NjiuRCTybgPCGEUaMiFk4if9i3xDc9m70k5u+ZU/+Lh0brwTQHKX4iScJ
+Z1XSBHgOp02P7d7Rg3SThA4u92/d/o2MvG+8EZ4R5jBjpN6SsZSU1cdkHyJ153vzgPuEXW4NxZr
wBsHFY5F6umqQZO9Xvt615jHYmJ2eg42ne8FOt0HxnhpL3MPLRFAT8mlp96Jd8uebRL+FQvLJTA/
Aoclclpbuwma4uNm7KbYVTRoYXunmsjEYpU42e8Cj21nEmea7W+/HFDSDc9fTOwHiV8eVzkIrwm4
0NlcRW0uZ8Ouj1+ghQnp3fKCOdFotQxEwuf/Cd34jON5mvXOZwNxPjI5dtfsrpe5lLvUjwgnPHWO
/XngbCjsMU4rYDejFo1Re9wZnJ44pG6K0nnQupf9QPt7mhlxGpE4ifBJoi8rpBPJtkKD7612V8dw
Y6xYNm2i5OCeLG0s8Xtw3Q1dCJPWntJPbDbPBBrenOsQO0ZISHtl9avrWr25qQxKuSkSevJ2RdMK
NAkpPBgV8hHVVG1EaPoqD8vGo5Su7wog6oY7sRMbkxoIcZnsyQJXTrkUt19raRAxklLfp/2HjmSf
Pvj07vHHyBO1ddRk74/9vWjjXA7a/ca+d0e0NOPIHQ+l1Bgdfu2pdgTv3mu6fuT9xczZYf3MHluG
jUKNLB7isPJPeCv+y36LgpWVJ7HqQ4K91/NJvWt5T/M7fOr5MBvP+lD0NW3cYN8C7672Lzxn6Mij
vDXehkqTTJmZSSVkvdII2ZvCpTNL/0KkW3XJleSY8UwyrbO6qaP4nDmxKlrln+Qymv0uwynB9JqY
t5R4A9S5vIogtBn0npMDIew3UyrfPV0+cnIU521ht5fVr/mHVNTQaV1ieGO36Rqdkv3rhFb7tVDk
KoTByxDduMgTtlnEf/1NVkzltJLEFtnc43cl/B6kXeF5sFDSlLQt/Auo1WkTKWhPOoEDtn9LRzEY
Y6UmSNBZlx6XD959XGG34PvyHsI7MXoMWDVphKjrobmMVaNgpydLct1ZUqAIPCNfLU7eXS5Mu8vv
4q7v9k7A+SbAAxu71nWdN+MaWIIfV5TN+PxCv8NvdMYr+m2iUcGr8fIVJCAlag3a8BzUXeupMJ80
FYEpeUQKZeLSlsAii0i1BukNqbedCPoFvI+HDaOFn8i1YoEvSICN7pBBhsCdv2RT3p3U91OI1jrI
1ElclBkZdpuB6tnJjLcRLDWjrWpeKAJXW7fVCBBSU5keWSFONVCefUWrYdN8LgXjt/d6JyukSMUP
nL4CK76U3lkvbZT7cSOQ6Qo4E/QlPd7CgaP5BC4bddQqnQWoSeakzO0WOW1AtqGThEjDRS4utMep
cgB/37GcqeKmVqOVzKpXEVAv8XEPNzOQrzFlJnf+KF9PBnaAlW1Jr0Poqdzb9QN+VLXFcJuF0i8N
UEwKuTgQJBpQG1Tv9QhUA/TCNsSK5GRGnhxW/dRLXZ1vFqh/HvCIQCyeHgxGia9svlnBF5UP5RyU
CMz8BCyfqC17JmpVEoSjXHCvWzh6+4sHDHWVDQETrLNi0IgWran1TJvsNiSu99u0P4RXC911TJvv
ekmkIid9Ybs4Io6dpPbiAIs39ERtWpdeuxpIBgqgVabuiR66kUbGn6KI5JZGju/F0Z9xnHahG9Px
zFCnuU4w9vW6e3WKDQ4huALN7SFEVuH+gJ1HKv7P82FpEL3DcJseA9PnTkCGWa98OPH2QtADVWVu
G6xoXB9sNlND6ZRI0qNfA9uIBmV2kVezM4zfBragRfyNbMSeWMV3V03S2AZm9yNXdPrQZ+qHRWVu
GNjEo0v2K9l+BJTTsPmXkVqljXMf79wxhTZbNweKei38TWaY2Brk3Nna0bGfChK9HTcRqgm353XI
u8IMbb1AG0ez0xC4erJMhYrrkMNqzM8wkE8FMBNcRPhGd0UlPAhjEXXYBQtGZKnlfiK/PQfiKTqN
3LwDHNcf557WCPSps/7P1K3kw8F7h4E0Zi+cN1tDhmmyD2g33bSASc/ZyLS9/Yla9kBNzviq5qYR
CPjxp0f1KhLQou9XztrQwQBCJdsNSWwVBX67VJiayRVNG39fBdsRqj6FTBFEPDGmxkMvWxsOie0t
JHQPklTUKS0E1XeP7CuVE58QNvLa3czV1aEYG8iIe0gFUc4vh0VnGybH9uWmsAZ0m5fww+CCbfbC
9p07V6q6VFfwYyE0AXL7D+rgWprpI3ENDNwxFO/sj1g4lIDZRpdQ3Cea0WdNLkFZWkFo42fnTK/D
cgEUNOi1+ITZWItcE0Bnwbb/zWK7U+eLtg6bb2MrkxMF+BZO8EzvxgmOxmETVUat4x0KygjPEHJt
thxmhkmIZla0JcmDqRwHi7mTYA0qYYYBukIJ9wV3fPiKMgMs2+r1ctoX+wSvz7Yy+OSqT5HGbhDu
Rrv2/4j/3v0inS4D6XMoQpVuiEMUN4EFCA4hCpptuMx5g9wBYxBEiidnMjjsizdZBn/b9lNIZMWT
KFzOdwJvuf4pkjiehuDedNEMh5si9GgmCWu9suXLmey7+TD13KfsZ8U9MD3ebtqVGpbjBfHIqo/X
bH7S09786/r7SzScxy+eKXPSx25Y88w4k8V6b8l3X44n6oSz+H8FF6lWZgl0fklt68xSWCQzR0vf
sJO4UwRzRscgfToB5t0JVbOSbSGx414e7XFsRg5iXmRB2YNlZ7pKWvH6hkNN4Dstlis7KJ5+e71i
pf1cMZOKVDdksqvM2k3PHAMxZAqJVwSFrhQpUaDAYQLS5DuRHV68AC/sb1MOj6Gjtn68jto3hbuM
/XTey+NB+xXCH+ZS87Mlw3+OWfZtM4vVWyUu1BtR8NpcUvzDJorJcT1Y7gV+ifDO3irRwmtwStut
+WWGoC2Fhb5DHizFPSBEZWq6kvO44WdZACgb0/X/qjkPYiu7g0n/G/h56EID+woUvRpOCF31Zfju
V5SJosXAKwG/8bFSB6wUL+hgkD4lRmjt28jcC5/FzczXZlkuBJ0WcE1lkXCE6O0bFE5XjIZBhVGB
Es+Zy53whg02A7X0onGgLrc2J5jEQ/V5pKCJCblt4Z/GhZBA7InWHxZ58pNPooHhos6mUhu+3BeH
0uJCXGR08i6Xhttf2XhzEcniq3w5zYdG9JjupMS7/KqHwK3rKdBdL5/HaUocUD4H9RyI7+R+G3Uo
6GCqFsDJPOyZtR1DR+k44BN++ujykqZB4h7YzD50gJc2pjNRdDEeHKABOflSPPQ7KId18/egCILR
g4oOL5uBkt0wGCHN7Rvm88pOHOdtDmug86i7810LBQgdyTFXYn9gM0FTL4oV9sHAzyr1kn9tJC6r
Af+pFxkpzgYpdRLLerb6WjULJ6cpw5u2t1QRZBeZVQWfYVo4xobumF7iTdNLoSpRPb0S9XqPKYss
CXQXTBhnm/B/3riRNdmT3JSs8lqlnqS83wzCqvIUE1LRuU84Pq3sDVv/8Q2HS36sm6BUVA9doCkf
ICJV3RlJ7KTMYoyJU9Yog7OoCGe2jtUh0fYRKzrD9pxAlDOsu3k09UQjcaYt9aDCnrQNXoDoBn/p
w7wdGfkyqSAQh63tGhYGUedcr2ZBy3NCN4lJGQe0fXbPyr3tW3HHdEOt3EKVGbNSO3MzpIbESqJS
LXZAS9eOJECR6dQcW4Owwtf1zcglxZmlAqOcnrP1LaXTXjfuulw/QN/FwxL2RFvyU0XOL6h/0Gkq
1AhaOeYLb96MEuVbjAfmQ9IVxgQuzRtA4AR3EHqLrXl7g/p/GRRm9DTQwIZm5M69a+KS+IQ53H8n
G6Lr+xYUvz/u5tMkSIMdoZ7Pg/tnM/LLWY1hRGl7iOJfqtVw4EUNmn2HW0D8miyGg0XhwV48Pyn/
K+NU3j2m3k42MB3oRfQUynMpHo9jaa6AxChQ3gP24i9k/i8TChw6kqadM/z/Fj2+pWgHxg1QYBwm
vde9/7ZhGhx9hDB5DekVkKp2RN+BXyWm7nYFMpFzHH+Oy9D7HBGXzHy4Wln4KpM1kns1gmNuT01T
X62m106o+JaZjz6u9aSisSjnJ5qeNJ3b4s5GGrlPF1rLgdZbLinSo9bvzNP3j1ABKRsiIBtjld6J
mPdGW69lRUTKEe2dxjvdnpENyGlDST3yrPb9wwVSrJFSzD1MdJgNggwDh0p/asUB/ffb9J7MQO9N
GNfkLpBVSbIT5+dqODVWT/fpCTNQcGcWkogQx4qE2iBcKO/meBfwzOKGDQ5diShXc8pJ53SM/8Lj
v4LDu6uINpiSnjFBCDmRY46+5VikdfcHpldq7g2BflX62u4ikLd8jrqXgiShcil5EKtF19jbGWtj
bs525901uKHZblQEjvfWvFDGpbLJk2cu6Y/Ij/UWBfMdRoJnrgqQCS/6zWajOTH8mRnOLyWHpkbS
3PmRYL4dncVAsn5FxbWpeXMzJyURMAfkQMMoMV00ucqznjs37aNxlQV24k1Rf7erSOuyD6RsUDRM
Vj3SVFMeYP7vSl0z51qq4DoJfROAq257K+L4PM7jTPMCwOxXjL7a2g/kQtYunZBL5lxZ3+D9htOr
YJxe4ILXs9SOqSZEeb/wvfml9RALEolqj9sYVWmRv7dAyTEP+IsEqmgTg5D1sZ+2gRYHkj+/4j5S
No6DNA8xLvFzYmu9GONXo2mkt+/bm7ik4kielVk60d4edP00yj/jWM+e5Cre4ZeW1IaNoUPvffYO
eB7rQcQ7s8C4Bbx+8BhFLtSBGaCgwWCSTlYGs6LK3H6pY7mcs7d99OmZVnv9MYlfEwhw28oUQS7d
feXIjHIX26hoBCmBvJkipNyPl8/dD/VA1HedNJUeHLTJTnAcvmitPGxLH7GOVN+TlU9HGfXRPX1R
zkIGU20+RJQ4z3RqcayvBmJYORHLW02w7d2qwbt9gMj3XpkZyIGQ/EAxAFEQgO2OKrtqoab5z6sP
t5W4k8TYYhMj9xScCSXgAl1JpYcd6/P3NzKQN4s46UnCMZxRtmeEu/7z36pJYwMhCETUlmweTXSy
0x4TxMPsTl3ThtGkC3fOPvVa4s0nWBHCKffKm0bLppF1g73OYgP7xYP/ccCpqVQ/Z0XA74BfzVmZ
yPNQt6jJb77k0myc5CYfI7v82FSKcZWhfbGSPcsabg6P4NKRiWE2vmKLxg4rWim4amNT5xl3MdR2
D17BLwpCA2HShg4xK6Q2KGXeYrRcrtcC0WkFKav2C9wME36KebTnrGfJ3LIzScfgRWcd5FKYvqzd
dgypgfi+9MGO0YjlVSnrgA6Vpn5K1gRO4NVQd+BH+sWjwXsFo2TtIdjBcUtWsgRdxaJMThyzQA1i
926pfnFXHrLclEMhHvEaOiCAhEV7/2gab9/YPTDfHOXsemP3NBy1uqNM2Im0X26bOLL7SMCu9/TO
C8n7YNOg5yJmFOY3XmwULD78aA/Ri4MYbh4IPrF9Y8wyEKT5y3Rqru4q5FG4s7uYktFGah3h3z5o
PTSHh+u3OKB4wjvxiY741YyCMBnZOpFl9gzUNjKioNGsF2ZnGwFdbCoyGZUsaT6zDEkxQQ82Bhbq
gbrNsmA0/kzhWK/ClBfLm/9uVWLZ5gilk4wpKG2rl/vBMLp8rxr/NzdhoNf8fgG7CdxG4HZFjARd
CQax3M/1dX+1vjSivg+/BS3T4g7frovuwudYhNMgndRP2Oal0wurZIHIpTUYFaZCKxQ/t4jBZ2RU
C2tuDX/Bzs1NB4uQw8M9T1a15M2ZEB9UNRKE1zEC7Dg2T/pQpJXseMt95ahoOlxKTqMG9FO53EnG
9FleT6r/eqDGI6eRznkq0XvyTKWiM8ASfBdKsmAf9WUpAxMvMFQ1tnpFMDoeOyMms927dh5Ogzoy
GLcF5XTsf9M8r6qWNexw/PW0VzTi2UDlwwzsUFLfaryFR4gdEBafdwdk7N45hY3B0WZvHhoWlMRl
fugSrorHw4qtuvxqtio0vsgjDUX7Ob1/fFka64zwhZqwvN4X8cAh/roK50yauJmJmkCpbOlI6KSe
/6DWMBiOyGI1sUPo1NF+m1nFhVF0flAU+rtU36qFWsEn5uXTxtN8gg6P15zL/rmA8esZ6BJA543I
lyMHzoEz6Cmi9APumMLp8aXMgfvQgcU5iLy+bGKjRl6QK5cYKM8CWFC2gphmvB/Hy82JIweSdwZX
j30EdMhx/onP6mMSACWNd86aaslzOHqT/W+toCg49+f6owq46NKW2pIlJd/cSP3Y0hXOKAPAX7AA
vQpJGDkvt/AZYQoL79a2JIHO3F1398B0teIBERF5fxlZptBFGvgkbUKkTqz5ellEdiktea3evRMT
SzoJQuoKJeRbrv+xmoPC0h9bn86h2HQIuj6+uZkds0VLM2/BfjSwFBvqEiX9jnNvw8WOTjFafnUE
NBt6UMh5FGyYFThaLg/h+LNsEvMfEA/JDDU8r4AWERP5akn7zu9L0YGVnJ3ceWJJM6PpvolikN8I
DfT+/3gGju2vy+TC0SLTPZORKgMcc2DW2aKjt2yCCJEl+htJgq4bRtLIGvEI9y5lmQaNnXzt5BkC
hgQdRie08CrhQF7rpxEU/Y0fa106scOBl9QXu/eKP1ZtSgVImXaknkUWOm77xxQN+E6Pow+MDRdi
JEuU9LRHLmC+3HxEmrolXlqW5ajNB1Jen7iClNYPfx9Y3N29uyTppGp9FO8zCLhm3/zUAHctMlc4
xbChnI8Xwa9DT+sq+cCbG4hF1eHMwbr4R+TbgP2ezuvXgsWSEa61sKYXlbUWPxzvEghbGZMdcqOy
Ouedu/YXt/a3u1DW4/TplfZGt6rwxIm6ZwmYFCF6dMMAGENiSy7rEFZeuZ4/Aro26LKAYVBRwU8u
Srqox0HBS6SUXIEibvYM9LLUGDJIZUMtmunpsqaWYsfbiO3LqbQmrrXZs/stn7zC/I0rwrAjR7DX
6Jm64mCI73D54m3K1Ky9ovqtWilx1Pv3shmDqNcKET9uc7D/04x0tvGWAiVoZRylFTbrMvatdyf5
Y6dRlhX+0UEotPEWiqBWrsTKrBsKg/KxUCYY9QpN52r3WaLywWngmBOlag2WIvAlahcD5r+1+oey
ZMETIFGEEXTJkCh1RVtwu2Vx1nnqsXW6Nx2IrJE3hcSx0nKlk29Y4TjSrrdeMvrERvHOX/KagEav
L8wZB28N1aO5Bp5cQ9bWzP67hrGFwlJPqpKsyiPqlUHYEqjVqOFqVSRsuP10fL9yXY1yjVoQG6mS
2FnX6VP8WBaav+qLVWzy3H4x6uNE1iUTEHN+ut9h9MGHGvwtRPO3O8MCSW/MtbSsKrr5+rvStshf
KjMhWZh4vsumih4CYCdFKNAUioQBD5yaEvVqtCienyRlZu9lgleWeynzlSF3uSnSC5opDkI0M/N5
KkCsCe3BtZaSgn6zGFz+p92lOyyq30I7bYfD14Z4GVjeq3ltyNLpFtMuzp9lPiFlTwmJ5WvXyJxI
z7Xh+BbyGPkrOU4Mfud8NPxsNR4VvhRkDWbo7km4ZiPThBnguM97lbqcTrrAbrT9RdXmGPnlep1F
1eR4EkwcXWVV9C8HZzij1xIi+P+QUSbflB4XeR4/QtDJ26cwENUnIYhTaeFJ9HXUiIxAGj+EiONe
yo8JogX67b5QM0AEicsmeBmfE6muSICTUjGfuo3VLRDDmVO7f8hbipGraXn+Gm7yaFy6KPz57iqH
By2yXcgySDNYdmmELD7aOSgjN+0Ki0UYF8kpz0yibTeuLDjycPCEJtDj7cPF1ecTSuxjxb2kB6/S
/qmLcU0kKoqo1kB8nWg9XSOyrMkhtks3fd7fFhjVsewJpsznpjsug1E2BlU0wHceNffn/hM0S/Ge
fTSsjNtE0p2VqHysFmdjUYZ/+lqhaV9PH/1diEiReRMSdkeckkyvoLPBQRr4iJcPvlwUCtjPTD/H
QVy7LU6hQptGHOsIOcOn3Db7LXLEhc8o5dl1jwtkkyBzq1uk15ARI/jxyq7eOFNylS5WO2JWW2h3
Id2bUNp7pJYqpskfcm6x3kPDIqmUevlUw6ffzpX1TcRk9KbejQb7bkcU41pL3MHHxc2tDhIAfnqK
lESNBaguodOxVsolfvTfeF8z9aAdw1pDgzxGd+GIsLvv6O/G52NSOqkcUi39fDV4ANmufve953rG
IPvkzpp5OXgzT8QOWNvVasHlSRf7PPMBdyrxT5JLrN4xqvToSPSv+77CelbCqs++eQTkj9xgHaBf
1pcLCLg5nANl+jQaa4r1eEuDLmIaOPTIi0S39HJIvAPn5IrVAm342v195swDvwJEuIb56GtNJFh4
jUbcB9P71ACInhiOsuRa/o4MSD6c5FH2oef7Pyb9OYkatQkwabAxO7s4etIWlGsVeyC7I4/MyP8+
QRqhO4jTTsdL38dfxImGLgJHC0wyidZ9AWeTzHoWI7LEalIOxUxpmkePCqPXwvOek2JigIfpue48
ckXXiFm7D6O1QVR4WnXkOt1HfMTIDJ61tg/idyHNk5WJVG1J3SzDCNQs0bIXZ+/joeIeZhECjTAB
+9LsckMBP04HD0Mh0xdUHf5aBB46XWYNrThudpN0QObyKZmU1LMrHkmv3D1MLmXGikNYtp5pmV0z
wzWsAGvIFVJnqXnVjRlA7KHWKLm9jOy1t73mXymkAVkkCGGsTdRzDHg2D5Q3vHU/HmAIY7q6ZeMr
jZvq+2NhHTQG2Y3frYYHgIYuwn2zCTB2kQati/5kV/GjqMZwf0PBNPqjWj5dH8NtcOOaPKFYxpqQ
XFS5fRTSSM+WYR7R6ZOEF52Vv9gG0EWcGO/pQegNE9DkCsqrz467gzMr1DGq9g8hBrUfGYpIqkzt
25pDd+jw9Av80IPc6oOvN9I3VHocVVmUDMt+jX3cII3devMZvX3sqKPHz1/lXLji0yhQ5TtkmiAS
9HBBaOGR6G8uGo5dG0j5dOXfLbAwua7+stnBqX9AtQyoW3iQb7Byc0NcEw5EEbe17qGvLXu16A3X
YZhrbnC8qrMKJVgaiaX8vj0fzDGRB8hMEDBm9M458VQ02P+KCCmoQMdiEiU7Rkg0WZhFH8Ipk4WE
Bk7x/QZzOsrFPmlhWph3F6APrQ+PjC7dn8gC9P3/PT8lkuCAVJbJ4+6DK/S9rC6VMgBGOPEPL1wa
fcibeNgXCWT9n/GSVBLq0N1FLedvyfV2OybKmvkSxOwQZwYXLKujxUoRhmDUKNdJU/j0LLLuOojc
nYDPGJmDDeLUKd+OFxUhRstWCaY9gpyHVfP52JDNiw8eOxQ0boWgZPX9F4mYdVpfLut9bUcSggMl
u6j9DniZahBcUT2L86hiM5UdEhGe2qMo+WtG5Il9O8rmEE1yfNLV/r1Aa3M7veAL4GOLh95a4Q2s
EiHBGt03wtpc6z9Ar1AOMd5T7tI39iW4wwYbRg7VvQQFhvd22vp1JNUrofWQOg4hED2Tl0llk9jp
PbQCMNAocdx8eToArPr0ga+9FjrkXr4JRH/xopt5KSUUYspyT2SOemYH0tt8lMOABBQEl+yMgTRv
B3EP/+c5vIRIwBTTnu4FTV0TltTYlmWyCMxChXFZf1HCSXsZp542x3+p+uC9rbPGOm68jzCiIbt1
BDi6LNXrsczkeQzAl+J83sUN/aPZVm712ggeJf8Xn5OXkcjs0mNN9zs/q3oaiDkvpa6yYcdEIkTb
erA73h7u9bk6fqNs1ntTQ9qUxJtl4qcX0ukRyfwmgW8gAfLXu3nJZjqE5PdIIQAudCImt7EEm3nR
6PWCZvBOuB9QwC3G30bpaMHLTqIcibZL5xZyFfEYb1HRWD9MKk0mVZIjNjhMLde3ss6G71khRBNw
kx7D1bBi9BXmDfOW9dGAC1/0qBmCHhq/FXsxrXloEOmVxNW7Ds4m78yWKDulN2/rKdeEPtAKHQGh
Fu9608eUS0ysLOBUvz5Cv/lJoSVW+nWdX8o9+VabJVPIEs6bKEsumvjRxVTJdioAJBfCCplLIn80
ZORSIwZIocE5fw2ZNdCp3LwqdYojlBYC9BUASuAoEjIu/HTmYJuXZc5fmFL4E7xYTaWPrmMj3pCP
XN4ZnOcOw0bFwhCRlMzUUHUFDjiLv8vZIxza39Y66XVXDKATLPZ0VSTCxp0N032pWEaLqrOJLQSA
b6/nnQw4bjD5J/prMdDjYfPX8iEIhYLMSkzuBSN1SMq8YXwRcOyv2w2KKACZFPHBYGp041NqxZvR
wvdMiXDc32Jl28iPhvX1cMqt70KN9IOfvHJdZtEdlTGZdMIXoAWpGxxAaQIYqPjbZBrR8IXz1tke
BkWnw5im2ppk+oPSi2IZFQoBF8MXBJKklpXT/XTPzaJgOzwWOxfuvsanvJXYnPH2OTbEW30jQBj+
R0J5QjKUiJ72lGw/VNMj4NdUcMq6RS9bleOVjB0uNKcT88gX+mAgrDLfGU/gtfps2uoejVDYGD1I
NIYFHTMrA0lZh+JdQSBzQqYmXAQhTxGSy2aVTljmTKRiwWUYVHKNrip5GdwUxH/ptLMfvP/84u1V
3XqDzx1mFUqUk5iTiS+/DvEV4EGfGXh6BHah0bWl7CEwqsv0dqBvRXnD4/9cJO44ewTYzTlyIkl0
gNX7wDG8UYMYhPays8Glog5o0bCjmweGjLGvh9pDgRVH/I0WOWJpl1g3ZRlgn/pZQpG1MTh9KjAK
BH+4e/uFuYJtOvx/g49PUShVIl3/UfyT0mnSE89sY91IYUKoq15kopDbRsrFunRq4oSFDbrjwSUF
/YKJjRwbYTRx7LPz+kNfO/mEmZpR2EkAYicSIAcmXJpSl/AJuBLzvAlRtFC3C0uXrEUobWF9qO/y
kvntspahRuCfYpZ8zgPc7mECwPvUDh19odDm+Yt05bZcBu4fIBF76FvFh9n70MNSzK06tffgHpF1
6/T+C0/G0azT7xqLB5ZMd1EUrO2oe/REfxrvbu8Q1ZPheA/lS6/JAekl8gIO5sF7VAZJS/ISKHpA
l6WskSCnF1jAvcWGHHWmQNlyxa5TDY6AHkLIi6ATrwPyVrI7q+Hxje1N1KkDoCBzzHr6lw/dIgA+
EKoZYJpD1PK55/VcEA8nSnqascywJiMRr0kjMWUoYzhBUF+22clhc2gl18m9MHleuWhrZMf5GEWB
3uo5BIPW8+9zKAPEDy1FB/KOw3mRbnmVNCVr0WrAN5V04Z3jTXQoqFENMklyFsXdfGY2wXoPWLAl
/JE1S3oiCJsVsTjihEoOY++g1Kkgg6p7rAAsmB7qFI8uNglhHtpMTI6n/6CvyKGR6tD7xigsFWmS
pue0P0szRYSGa2+9BytRo8gMibKX6pw9W5k1larjot78ucx0eLt6DCeaEeblolSmIlUMeGoowlYn
v/vLSz1Y8LzPnNsREIln1BFmQl8phPgLNldC/VEdH4GPIMh9JxvmmaOS9TpPFUc6mDW5iDf0o+Wy
vnmJBL58zOnc6BGBvx51dxrVmgsdS6yH6zCNjUEva6WxJGrD6xEuyKFA7qWrL2bTQ+sJzY6gwuTM
997wCwEGZeBLd4sP1Xz3DEArvIwGkvclZV86XHEL6qV1rkGt3MFEUVKB3jwNOXblbwFEdz+Zm3wW
OxkLPurp5NbFTKXcmU/gwF3yAGFDevzU8MeNAxbukMA137o+YWhbxaHxt9wc+LCzeFj63LvM0d5a
Q6G/ZHe03FVkHNk4/B8qTdPhcE13IbBi3p26P4a5ECUnY3h0nEzWEY7a5eWpx6m/jOeUSPgaXlSj
xUrIroMvsEqoEE8RFmZUbFYWCs4Cr4fzZ/QrfWLq/PZeBpUilQsLaHCMVjY5P+pc/N9Fr1TMB+Ga
F0FBGG9d2w4YBlEVwOHhhzfvpu2G4F5KIrjw64e48Cy9REl9JLpX4Mo7tJsWE+urz/O0Io+rrPeC
AcyHJnzfI6vS/V7/OAA9EYR0cfATDwB3HXn5XDVZ+4iDV601km9JHlaqutFducFdm1BxDFJBrdU1
98oQc09W7TNf9Z7/yxxeRq7+wm9n/1nBaC2SCATYF8J+qnG9kllQkmDF4ncM1ku8/pov/fkkHZZK
GU4rx2CyHrZASShIJOj6xeG4CrK4npChqmiMdLJN9JjmDh233vn4HwNLU1HTzaC7JDuCz/K+Nmu/
PaMKzhCjQFYgDWi11D/+POyL67U5KZ4yaQCJfaCxbv1kbzTIjJBSjiq0wD87Dr/gSr3kHVjCzybJ
v7LaWs4d26YnmiotzdQX8e/rU3dxdZr9a/wZ1085bKxC5pSDBFhZQ3I4uhS6epVAxDOBijk3+SxK
t5MUV+9fOTOex7eZk6ICuc+8rwZT7qlATjI679XZB/yKiLWVQxMPfMbXMolokthnPugz+yT+/pf3
+YqcNh3I0uXAis4HEvQJ4GaemB1leJmQXOqqa6vWe8C385aRhrtyx2tGI66vs370iCPrgYYBy17f
CWu+oApu8AjjC6iT6rsqrK0Zq3ocbY1KJyP+V9imUDejMXiLQHwx1EnHc3zfE12q5lIXJv56nyvi
A3KqemlMIE3cbUAHXQniAH41tMyT3XZc/XVZP2SAyb6P3M2dMBqpv0R4QOwDDyAcaie9o9CVqTSe
V9QZrRNpNC5+nFEcGfKlE0rdYoUcLPX8Y0UJl/Zioqvx/BN3xytyQYG2fKOFOcsUlzz91JQzB+K/
yT12Rs2GiFAUfic6LVmb1xXrguuU7QxF++TmvvIPrSisD+k6YdrsSe6yRGVXMnppLwCmmuo0Bwuj
GAxvWktLfUtTKogJMy1EefUrhkCt6/6YBFZEWTS8Rqhyp+SI8poy4aI6e0FFG5vWAC3xqyQbZPC/
MejvgrkiCh1J10zOC07MD0I/rTIKiV1EmcjbdkSq+9xAbJ8pJRgFt8xY5/67PjEQ4jr1Qwd1+L2c
o+11JUa96oA576Dthtadg1zqBkRL5K/Uow2EUYCdvBHG0NMjWhq+vJD7lWZByUeL4nCVeXzrtUPP
FHHqa6GvuuYsLGeCN8Okl58SAzY5VclivkT7cO4VbesuYuGUL7Pac69TxtYPLrZIpfQlUuhSoa/y
03tmqpMw2SUuiInEtIRnELEe0Wri9Z7tYsNKGbQuEfQVXfc5boSYJUCUgFWMiMD58R0DEWzENODX
xlG+zPv2Hols1O7+JP3eQfxwECNX8npvvR7BZD/5ws7VXRVSifeFjJUqoii901qtKd2A9ZM+0uH+
jymqX/+IHSX+IgeC+eZAYtLfVShZGie/JkcTf/+upv/PiNrCD8IZz4UtVEtdf/mFRFl56fpvFPsz
8VmOzPEoteUQW6jOH1T2Jx44APIhjFG2wuCWFnXnVJ7EChgOhJLYEGCTHrGCUxPeKG+7h8ogIDYU
m2q9oKtHbpnXyHEHCgcgpH0fI0NotaRxzmgjMgPFDRLA+GboekX26HIXcobwQRLedQwjZbi2kePv
/XNSY8/lLnn3g71JkvRkPj6MjcNMLIyPIGGFXdvjZwQDBYrSfNJ4SZiN6rRZ32+0DHXYKB6OJ3U/
gQ/Dy5hnZrZgp0juzGwXMszHIiZNeVBM3KHz6VvRMVlZE8DTrzmNfy4p1Aw/LiTM+dToYe/YntG6
ilZ3q5+wt81sjvWTNd9OECbv1wTdEHrykkOJY/NHYuQNyUI+Cxkm5EbC4ADa1+k9bMxKi0WhPQWl
N6Q7RprgtzKcM+qZnvxjVUGa7IFSKdvtSzINCg2BAXzDpd0oKt7KzBGzCVIobg/fLsDmhskgITxH
cdNXXWxlFKo1q+EFfbqLIpO+eQb23vwcVimkCPRg+ajAJReax7Gj8RvPpx1ljiQEFnWRtzr07L7y
9GqVxaniMFNQOCbOIKWz1Rjjt7R3j+cPyR2+9yjVxpO34XW2kunff1w9IvrGxkoJYarnIie/DD9c
o5kk8cB9xaIv+92xdjrsoVxN5RM+AVo2CxZRqNa7IWQ8RGFOBH5OLX1BJ9ZH1oKFI8ImiJ67oK95
tS2DkY69sVK0moqWXmK/B6pNCBl8qXlpexEvvWYeRZdOBWKV+8LZW5XlsUFq36TezQc2T+9qyITw
ozOntt4cfFGTCfBBHNvPW1wP9EB2+vo4qFeH058ZtAZ9LzThsk3UC3lq6Pr09v6vR7Pq6DuJqtNF
vpqFAhYodFkG6jVCas93n2PPbXqLDu3WW9yWS67smJFS5jJEa6wN+GY7r5HmXiQ8d1ZxOntO8D8c
mfmINsKhMwHp5Si+UlYG2kZsu8EYaJ+odzJBRtgtWYroYyjp+YrkwSrBpcWvLOTW0GtnfhTs4Icc
ARr6Yv8TeYfQc468EKZUIpNhAZeZ+tpJa2BctFPpVBFQ8fYnaYjmV/lEbBNjq8DSBoGSb+NNaHYJ
VkVKo+uVV/wnNb34D/i15LVmqkkFxyB433sR69HeJINtb/PqUpl/7hEziaxMxts0zWr3WLcv/K4l
VU2HfLZifSS+RgHS/WOVd7O/lyAh6mGVBwPTYETU/1c2accmETiPEH3he5dPzJXtqlBk8F5xYG93
0vk5DImdsp4YEIRwalxlM8C638VMa7t5fZZRd9UgYcQC4rf+c7EwoJ7WQK0vatswrxk312Fs0UBB
CuZ6pQDeix5NyWrGcO/kqy1QjHJ2piLudWzAmHMV8KGFKyB3hCZb47lAPTCG+ugL06CP13o8+iiy
RmGlDG4wPtTqG/nA5z+5JamOGgqj7NfHMlAccHNcLkQ+sRDuPQTkGOjshCypUt5Bf7lZDGjUTadv
+b5wS6eHEhTIEzIXsAqGpNjTdrDLmMxeLxhBl3WSgEi3X/xnV2G567NoA1wZzBJiijFo0B+0sSBf
ECqa3IbNqRiqPQK9pJKo+NbEyLknpRh0BcZKxEAmZSiDyo7sb9GhTiSz97CSX8RofwgHemaMe1Ww
O9wVJ1MlM9e0Ef9+6QDk/W9CDo3pV33VazWWzSy+L7zIXYblACmP3jssF6TKJJqTnDR8xLOWeQh8
pWgLShxyd1Dy8MGupgxVTKc5GFPXkXDILAmCCRFCkco16horySf5/iq/Au98VourW7LzQI4Geoiq
q/cBzLXKCt4QIP6zk+AvFHelGP/FrGjiGQ6KZ9FuaBhhuPBbBtc+0G2FlG9BcDoGnxoM/weEiMcd
IaP7hd7VT+uEMGF/QXehNZbfT55Sl7CM0SNaJ4XPDJsrSVCIvkhfxGRcemIvqswtzznynWApmlQE
P55n9cb3E0eKlnCrpVmf6WKQvaHCaNpUOMxo5bB+hV7kaoY80MbTp67ANMBuDFOORaY1b66BlFzG
+8c7+RZfCzXm5LHAHPoKicfzaUkxTNvLixHwKZMjAJ41LvKEsqRGDfCNj93qfiGCLOSPG4e9nMe0
PIbV5qBy3y/tFS+njcVbfQWwvOijjth2bEYZugWjso5LqoAhM9aohqUs1HLX10maS+WS2dhRYJQM
ntsW7aaVuAd8SOtxpsx3BdQBE40EH0fQElpJOB3tlL15IgPq4f7KJPPmYybs1KssnER4iQp8okZe
wYQkt2CTioNuaS1toXig9wTa3iZ5DKBRv6huQQv6NiYCEGUTvjio01bMBLjxRtrOddfEUiJOpjF3
6+cThwYPioPxSQLwp8f6kFxlsPfX6WqqT8xJMIi9y/vSzpYHjum8NnaObrJJv1XOubBah2Ot4fMh
cXfXzpWl9D1br3aJ0hurcVNUqOEvGrgKpijgsIp3uflwWbXJSDqaNW50JODSL8WvrnnvSxW+FFVl
DaXG+/AaE7xn2egkGN/HvlXCYlQ65HaV6vB/TQRUkZnbH/zrzXg+IjwIF+biE1kS51HiLtgun/Qu
eexO/SnxjLTcMdww+6v2wfL+jYU9SeQIPdenwLDmuzlbG9rEjOp4N7CVGhbeHU6mCGZ2Vk7NMkTl
5OdIJ4yolzsMwSKzf43IE5on/+rzAUC3Ydu5xTedli3/GB5xsFJhJYi+5KltX60RhAHILEMx3Mtd
gsQVdp8jvWjl1W43bYthf9BOlLQ4GfXUZkdUjIAK4/eB8eGd4UwKIu0Dy4VgIfexLnaZVCY1w32O
5XqvdM1PhIRMOwZs1haQwe1s2TYHtBFxITrZVoR/8qaKzhxJqBHAuQEL/uyVTqHkyMl3ofD6vZND
eRMzLcINSvXrcZ8NpeFjqOeE/04GHaH2st3wddTqcvl1eyaql7sDBLoYpNHArj0AJZUP6CeG8joJ
XOzQgfldb+nDPaHX95knDdFoJozyCZwRYqyVLcCONs3mQCzNGgjk/C3pzpyji30zNLcezPmhJU8z
YEwrgMLGN8isTx8Vc3zzqjwK9vH6Y26Fmt5WGbYTPEgicgF83uTth8Gi297q9k3/uXuz/+tptIcJ
OU0Aw9QMrRTxkzmOdQO/WivzKo25zvC7wwqK0Xi/WqyLwoeoWhYB5IubyiAr/pAmkPcyGH9fhOA5
1b8SHjBd6EgNwHgRigZavY9XI4Ob3YveyDpnA3FDwZePbAjKFm5azG8j5XeJAvoVbi6aArPwpt9J
WjbVuQuSpjN6S6KhOc+hObIphzNKLGQtIDWEMsAxBqYOcRQ/mC1UfhGA6zsFclhOAybODiYBrPFJ
7gY2haWxaUQbxs7WOsdRRsPOQah+BovA9QlrevqMByFW+A/B+pZzc1xazqiNbf4bX+dQpcDO+HCx
zW3Cuk2FDIOXprB57EPy9V9jLPCdlQZtgsPBVMx2ZD98FIg5bjqBSFHp9AHUr0D1ftEfQNpEl3uf
Exxgp0qBWNFBnQyHqI2CIYiX78V6HfqXXTwp/vnVGS22cVww0W3BEGMLT4ZnlLNQ2//Mm/6UHJaT
qKt9lOie/GludO8T2KzCz30Sx/EKG1uyDi7Uq1fNJLFiyIOS3x6CoFq/krYm8VTsfJcuNjnrHvwR
y1zFETKvaQ7EKhMG1srnXH4KLtVW9E92d6jEIQ6w/if7QKnrz2XqR7LAXffI2i5Ov8BBmeoOMj6/
XYKwmf6xTzxRft42qz87979e9A8ZpzPDmbmOwLEp+9v0D9BVtpcDljWLBo8wD2FHlROsA4dBz2Ye
LB52kmywgtAB2smk0hVuA3QbGH7hMuurRYJSseTl7uKaGDOR85tnIJvISCkiRPKRoGSZEXgMt9vU
8rXFgM8OqdYks28lfNg2dS/mGIIfyuA9bhZhwOR+RYeQr55A0gvGCoDA4u2fXBeDGtsu//EhHU+Q
HJwEib3+sCg8MYHRLAzuZLZcTbbi7mLzTz0SLwvNr5kDnn3AJtcDD00kehZH7xfa5KvOfjQ7WoX3
bDQFbR99rBEuXvSFOlkNub7uyEpVzKxUxliCRk1PNdYC/HakjdsWLxaMGH8OMd7zIgdb3tAWJlMP
CAZkjklkXMIeC9qzTQrrJ7nDjUO1T4hVUGsFp53qnvFzRLgjd/QdlNGOqxXNNMfmaOYu70x4Rvgf
tH64oJaDmcCdoycJkGMKxI5nnMJwgrvLktQKwVHZembGGwvJ5fMdyv4m0zc90YlzJB5oSlQgfqTy
+pdlxNJELMD4yY68WmyiEx+jc+rtgltvZyYPoW12gtek2xsNj6N7v5UZfVr3QyZYGsDHMVrNHDIY
8OyjKXYXOIV0xUspJnOp2KgAmZWFUb4sYBlXmA3ghFGcK+yQGM1yKKYfaLfnM4WJIuYzMktFoJ7Z
mIlJScQvfSkDqNGzflVc3IJ15u/wG4Ts3YfrionH4JlfcnLvGT9VTBB0UdSi7FZG86qzvaZbOFlh
YWE7Fj1cNsBTF0EuW3Sw4181jOa71J1A64s+OiDo5SOo9D4SOmUqgBg2TcPvU/SvYlqI/iyBXEZA
VCPSjRGgaZ8OfkGgJFfrlF2+8iuYy8rtbGc6nXeQ0tAoQ9R5yptxqVPrr0/GulQKX3tcbK+TIW7I
/8W5yo7URyWSZv4J9soJ31EexKlv8k82k2thkLOoBt/i8FVKsfIgVnSmZG+kJ2ZsJCsTEQmWNvS7
WdR6GRmeJ2GMsOeA/Mn/Jd0zNBQ0rNHSGkiQLG89+1PTMsNJY1IGybYr9+XLMGraOMQOI5r+/WYJ
3kh51FAKiLiCD8Q49AEAsC5qOuP6PhAKaetwnV7dpvWeVy0LR2SHPZDasZugS76Lql63XuwIFTHH
VldvbIBrFURkFfA0Ygl3RE7179hI79HWLOd5XXcmNSiqTxzCLHgQyv+iyGIyHx5TMLGXryvHSrYz
zjCkNL10VkDST4D13SZ6n7Sn+LDlb9vxpGDhaaDiry77GdxD+QUG4N91nGmVdwrUX7asjo5RB+R0
b8EWAUQMIJCMAlOGMu/lmNFYsPfZBBZzyONJV7Dkb6nx+sMX2NhS4oYSgOQmUHMaPBgHuGwkO9XD
tsG29+f/BPAutKLJfL/p6C0a8apLrhUcB12bZ9ptL2sFQvkqP1YF+Y4Vuuqn3EKgR8rpEqM7+/w9
NBnryYzLR0J4XcjaFLqOliTXi1XN8gCVfybUE+2WY8rF5ze7OcxKwFGgBBB/hrduko2Hv8GNrBSK
u5hV6jmiUyLHEJBV7PjiFs7tAi6oTo09pgKxrpPhbDKJ+UB48+bDlgtbG8+DDM3c1ICCetzLaz/L
3cgWO2vuTpjDNNO1N6cP6VG3sq6kXExC0kqArecJ9gQwTzyqDjfjghs+JHqCxyUhYgWKZqP/JtwR
jV8dTZIeoCUtADjiBJ3ky4PI8n6ig5Z9X6Jc26NZ3SWOOFaiB/7VdEqOrIgitulP+EVqrrTYDUcc
3zbHFmPZzrNOltHLhQFEEM/BBJue8yW43bnVzsl2UFPAXROmkJOfrNwxkDq3aXHW+iD7TL/Dm3kR
knhWp9mtBOJJ2Xjq4Z+dJYRUkx7Qbj1EkgDh2vW1yPzlIc4PDySXVa6KrQ4Wd5gg+Hxsf1fFQBHw
w3Mah4bUunXA2DbUL2ErpSGt3yWDKjPScVgBkGYBCpbHy7Nt066KsuRWMoMdyf5pNldc/99zsOPT
n8c3bL0l2hgm2nunU8V9Yv7r4Y6dCNvOf5438b+1ZPK5LP1szwCA5WbOYkJIwmpcZl6f/tLSNMb2
dpJcwE197zxzs6AeZWT6+gftwmPL7H2YOPjJl3CMo1oXhoQ8UaCLgsNjW0LhAbDnQPsonaMeYqLv
ufeiYVMN/RuLV5kkorGBKSz3+Xsd0JF0NFhnkhBY1TJ8vFcS5MDmx7ZPe/SpxK2BXBLbdqO2UzNE
+MktPpxH6ufsuIUKaPpqCALzjBBitgoUzXghogI9374hd34kc5MpQ55BVB0ndHUBzJEaDPlyAd9/
Mg8L30UyQaair0jr33UPXva9e5GohAbE5yf2T+psR2W5u1HBgtD4IXipdFZ/87MqbE6OEL2V1SUp
sP9LXqiLYzuZ6qvfATH3XhIY4ezlcM/1xRPvuZM9a2Hv6SfdZ8tDgmtX55x6ZTco+Ur0M1JojXs9
oM6vL/MTp0ITJ6MurnMeJ8dE/lPgF00gQ4DZr82lHOu/giaZ5BNpAmWtlIKLvuJYpQ78EkED7gzf
9vHkeh+GpTgOmYwIXpAQY4fIjmMjYalC6BsyabPLQt4NcIiK3gzss+3B34vONAhbJZnbO9Slhpjw
CEMOW+8cskX3QMD7g9nVpUuFa6/Yh1LflGon0TRUvnAD4P4sLFTNhiaJTN/BPtCDZkoVcwNLH68g
+dfiKgpR2NUhozXBSdjNQOVwOgGJBTOu60oUOMiQxV5FwO4ifrrGhT+1tMNQzEYUqaQRAiot8uYY
WbKwoC1kmr4Jfw5abiWfsnP3oEM/7kDAVP1qZ2LCgSYQIoLE2v+AYmkEQ8uLsfunVy2b1dZKtYDe
W6m4sIK8mI3qmPwW2552ox7E74Gpp9hNBiBv6dsCC0vYkE9JHJLIOIv17Bcf/gWIqTTozBQdklbm
mEmJaATn2H1h+5ceAWNPkc1AGeHxJ13LGxHytwZJ+rBI8hTtinDM3niSLjJzgPW0VI92csnWgUVj
AGytHHgRZ4vflrVdGob/OWXvOpvbcPlHuop+7bXFpg+YF5qsj4jVtNoWJQz97kqrNwEJ+p6s5zw1
XgHfGvuPvM4JaPg6iv1hCvKgssi/KR9tUS6i+1lxVmRfcI+NjN9mpmiXxGIxu53+/AfKIv2brbEO
Tuuvanp9OxviknTI0x5M4z42DHwNwa24D+C2yycEwM+IFf8EJsSF+dL1pCW6kbhZTV1tSrAEtmZ5
Rj5EgZfS4hroQ+8KpoOqa/dXTQ3ZUvdCHzQAOv/bmoWXU5QpoX0ZzaDRJ87lNmC7q5MR4s6RBND7
oWjBMawDumzuIaQl3k/D5B3x7Lp/g9i758LykWGTMojMN+5woYJU+RefqARNO6nk2Pu/4PrNe9JJ
DdiJSTgUnTc+7LKeatjkcWB7ngSdksTfdRpUpC/q7ZFjDf9U3SLYQNNy+xzuq4xWZwhzblBIrlcB
ZST9TVDvISmn+ZGRZMUAyzcZFFQDyECvtM1ilGkV/8Hh3WuEbLjQpv63qgv/J2Wx1y/EGXdltwZ6
EAOmAG0XHlChKSnYWW38mFyzAWji1Yr9+GA31ZGedgbkcwvaGFapxgAfhBmkCPeNFpNkLzuBUzMc
Ml/taCyBEQvLUKgwa2IVtufUxgb09jhM8iN2rNpZK3VTH8syuobgVT+YFKzioar7h4ZDGC3jbrHM
vN0ntFekbzS3cO6LTXbaEpsE0prctxafYX5PM6VZsuM+tts9e/666DkHWePBX1OpkO6S7HDnF6ds
DwoJzigJrna/3RwPuSreDO6LhiAH0For8vgFZcr6z5qdMUT/18TgFKj47BEIfr1yTzx6GuRwn2R6
1HUwhQaZq6dP5v6acFF30KmnN2juZWRAK5kkU60KZRJShgbyhxsFQYfvqyrYADjMJXxB3+S/+MzM
TpUX/c1NayYviPv5qTvzsiZLQoEnQhlT6twqHAI0SBExFlU7hX1W0pXHWdHDNOg4xznGSTJzOuFT
z0lgM8EiyamemAjfw38zfA4PO1RPhnDj6c7qpX3iurtUFvb7bzay0+MscWc0QBbZjXouaGjPqdly
wnmmCzsCFRbq3020HD25BUo4LowBRDQxzx769XqYPx0Qket/csMacs6VQ5QxEVDM2OfSfcilTXne
bfoRp+alyYGMv+HP8zc6/ehUnUalV2I9aU9giCrYWdUEmnV5MP8lLlZ9sNbu6aD+PhYjQdIWXn51
NQHPaGkOrLKCUz9Z/n61iiQOC0ySsvQb878HyKDdFfNsVWsBoitiRE4atSlx0LZvWOI8xSuRzkGE
N+86UzbgflpWUC61oPEjRn7OpVQ7as8fRZsOK02ZjPt91Ex/GThSzJqkNWRIUosoXYzk1yUZkAX7
PAXrMQKB/2VSZn373TvAEkYRZT4X3eJ1pcXOp8K9Fo629AUvUDaWaTHGWlwl8X08Bf4iXG/fQm7Q
gaxI/HCjpB30fYRiZFuFNf9kTT1fmR1A6JlZQRZ3TeR2yiIe2ei1qDURBXRNSmF7UsD1Y5G6JLFN
lrUOByuVonY4RoTfxTPgrFJSWanZuAq07c1VZZ2CB91qpKCnVbdmeKASXRNIVQId8Gi3E8BF514+
e19VltIXxgThisBG5/lQg2kOt1l2thkwofs1QioUILOUwAM/fRchCo7hWJC4YZw4tBzCKFTRcFTQ
zplIikOi4mymZWUZRWC3gRVBS4p468X2VbI7zoaf+2mWWyYndwVxoI30kXvl+EJTiWZt4w8VnULH
ppzGl5BiEXPEVCk0D886fuNskMJ3XIVaFYNlaDieDl3UXlobUcQWmfToGahLZpg6+LQ2lEbAdMGi
x1zBDrwPEhvbPBr26enG4i1wWAxMigRAsaY9FvDgLD2p7tnlLsO5SWRZgGHEYx8L1NkmCdJ/V1qt
wRGcj0xWNgiKtS5RYzplCPThF9zAyKFAixe9J6GPjW35dc2c4yVxaLQuRG9u2EAsYu26C4YkFYbH
GThLZ4KgGYWK4QaDT8Cgt5VVq4dQQAnXTbwboIxzkjOI7JQOsCOqYfctwRdXXDrx668jpi2f2OYZ
Xd4/lldu+tI7ryUusogqBW5qpR31tJazQTTqnF1gqpkCyR8nzC+/dqX+1gh3WPpkQnB1SabkcyL3
1mGgzVQ1XKJip9QOKM359aMOwoXttnAKKznRqGq8H1bbOhKoztJIbgEe2ay2iz4Xns9MM/2MmJkt
VnvdfiH0A9tFUUVF2EBktMtptyuZ2NRBxHW9JZEq1GcaKr7SKqLSv1uFTS4/gpZQl0MYIbA+3gSP
Sa7QDRW5MB9D+WZdxxDQVP7w/Msde9n+SA5MFXPS/tCFEFUtjbAtuUc2R4ibkuoixbHhqaWvi5O7
QudKycZL/vZaH/1KWLrYbRXQh0lSgSwf5QEoPl2F3Qqw3SUP8pSipRQQNTy51I53S3g8JLYzRFfs
UQ1+GVBH8SkDx1Jl5QZuxBE5du8AsIJAhL253SqyGO7Kv9wobMZPPYT1XVmI9c2GSjlmxGF9VlwB
XuaOC8xu50t3aU7/cdYMJ5IzZQk2RxxOD4OoWPIrvgE6D+0Xm929lFQBpidnI30rMszUJbx6eN/S
+gzKOgThtTLrOYvisFlv1II6FwjbTUhtqdQaQjL4GSsA7B8GVHXU7Evymyo5JnxQ6KiF0nW0S/yh
Ja+EvrYMrRK/BMxc+DBeiYeRiPwaNDUOMCCk4c6LJ56Wug9Mwd9urtdnhw9lTV0CbpbT3kPOhS9D
cK2WGnFfZHW1A9R4fF5ac39lpxz1yi89JgZKSxsmEEW/IRTc7eguvGoACkU8uqZiY4qelncpUyNJ
ErtVB5ybu+MtlfGLfxyZHbwA0Od3pkgLazKPJcIXfdiwbEGbQEgbOcEdtJeIlE16KfPVMJKsd+IH
1TOYYMU/4AsUerOmKcwtqf/kBF9IYurVD6ZMcFwwh/h5ZgvzwkMCW2xDxDJWjPtWXZkzmkKYS4Be
gXS8Ea4+TQCfUG3x4tWXIX2xxQP8kbBpHs7Afgef5yKGb5bugby/EuALbAmqPpn9PgGIsF31iYZN
MzmBkUCBHyNzvkzjLgT+ROF9KoERNxWw1GrBCM2OcwNrI2sScMBI7HoNqv+ySzSJeZWLxAFEZEP5
izenQfB0nmtPxnEcAjJ6W97J6Wn/4qiXMIijdT44H9Y3g7/PH8pt/A6WboA+VKu4Fz6rt+H005Gj
iYJQ+jjVmK3I47UQqHwoDKJkYTQdJkVjoWm97SkQdF9swJ3+Lk54JFDcRUAtrJ3/3+4zNtwFagIy
7XUEvBmSLevy9HrMvW8SpwFNQP1Abd3cEOZ/vF7zhJObgjITs2S0B+gXTKJRRwIGTLY2SFsyM2Xd
Y1JL/dmnP7DcZEPhUDbWmIlwcuwaceMUqVMicC8dAbz0D/uuY+vFgSOvCClFcZUVeyV84kY0uR1f
Ca82t/ZKQw87aaX3H4mKpU3v/yFqfwC3AwWUH6RtJGzCveHk8VXG/Z1/kBUnpmsZ5hecZYa6DwjU
Pt/xudz5khRSSNTp4UnXnif/EeGfUB14QcdcEvxW9e89qnT/At8pteHz0ougY+JSGr3zvm5I4CiW
Kyc0sI2jSk0Zxkrcl2dj9cygvvW/OvmFFLwqRmyACeTJq4owkQO/A5Zv3ARsvid/JSTeyimmpQIk
j4IMNElpzFSaN8baaWL7Pc3/b3vdnmj7eluq5yLJpaACkbMmUEj+L79cPDQU9IGMjeRQONnJK+LD
/ci/c5z3PnT8YewKfyKj5L8IGTDdl5AurXCMbw8fewZRApaRLylVoK5RZ44NEQEBzgVWtEszPMvC
8VpYGefK4MsVqmRZf2qI7ygZ3r/3W92fjGJ3RDtsWTLeoOl4vUmxf2CnOrVJIcBggbTuHcS5fJcX
MogMaVUuekgSp1H+X8SkO2eoOWg4gCmyoccQMO/khZj7z4ouKC66MU1L+R8cBO8R9GQJ6KnyhyZJ
hJoK5JAbXm5stfLCyfxmTdSIKx6p2NDUSSGuCjQUGjVBb9Va5N02rKY8wVm52fDtHpZAV1cvHkOp
QO7sxwevjThzLtByef7yn0L1VFJdXGLiOm+BMTjB/3gDdQwfX6Mtg2cHShRjusdJ3/vIVcIRRF4T
65YDrovIF0UlirZqO9ffm7fN7PsQd23BeFhTzurdYP/dospok4nX0cftPDYtJq9WXzt5dbZdQoiq
m7dMkWA2gqV5uivg0f0rrjIJh8pwvSGBVTpxEGMhx3YebJmOdZYNYaYtd6JRhSrY7oRS5Hdbnbf3
mqTp+42IZQTZBSQg1tKXhcmq6vBoYtfiZ/q2lxDhe/+kXsAY2d3QgDuv2x21hGJ3J9y2TtEHvq5C
v5rzJyWgQS6dmzGiOluQTgtnmQBYDqSQ/qGXWUpBusS8Zgcj5Zyln/4BUDYtCHXt1KzTWc8/ROEs
LlF/KvzE7fk5LKfLXpF7tZGbmC2wE1LruthuS1MnZiYqjIfdy6ZFhVSM15e3vbRupO5n+ukA7tdF
Gw7aQJVw0IVg7ryOYXk4ZdlKbgCsnsZxtKSgIRPLgU0xOyf0NQhPC87wy3gm+iAtYEZ7t1l+G+4h
NnUZdIFrvJjpWw+Hq+3u2NVzRcppaYslmxv6YAPMOFtN6KWw6IH50A7bhe1HyehD7Vodj31uLewY
NOeky2J2UPoOdXqcSof6iKCO3CojY99tanADw1qMt7icG8Qgjsge9xa+krOqAuh7jduE0YKZn4TW
Mvl/AOdnzO7eqkJS5EzviSHbXXBzGDlSI/C2CZNS7gI3T0Qmwot2NDPfI8B2O1aQHeVBURdSWJCu
g6TMC55wG467seDYn6Y39kRQ4j//4GO1qEmHxDkdOPZVpadfijet4ZngUdI6z4fQlKtKCX3swy71
2eiCzbncKkqiXcbQM8Nb+yS4y+jY9I/FtFCZdxMx1UlKAV0tfo9Ayq4m6XxcgiZtafKU6o31zib9
X6sFaBtEvCb0XRwI/hnOAZWZbxZTuxwgcN6VnBRYieSIkdB5lnOi/WK+oM5Z4mBW6V2aeW1en+Z3
xBaq4BvlGXv9pA5EFuYJSDka2JIWX3y59oSQegaMio/BN/JP3MoN2sYs2KlNzTsOyCaEOSFgLEuG
vfYlXVgenDlx2Iuco80IYmtjmuQuV3VNVhFvAp5yiL5eUnVSjxJSgB+CpSqzKBI7AuMNCgnZgHMg
VkNxfF5eYx14xKllaQmU3EDB+9etSmvw4cRQ/7Adl6tUE0qQbN/kkVQPr7fSp2zVqIn1GCXDt1Wl
RjCpkJTqVPsNfOfQlgeg0dpNPzE7pgzS4FQFXX0XjzsGMU+z5E9P9HCQmOF5GHgVdnSVs7vDsdFr
hLOJvLCpIfaj1p9pyw33+JowrqMT3pILXraMoJjdWU6BYbLckHRRrfoiqXn+8xfB28fGB2optHfA
bafl+4/xRyfSBien6Q9dI7wm7rqXqhHME38wU5rDJfSutOplvMfbKTtjefzDaLAaDgC2xsg4jeAW
4qWshqTnFGjxFLMm1xuYN02lYR463LezTg/OrDQiTSc4ewPb4VFo+M+6Mz7U3d/WXmMAyhjbEs2J
o0SDGY8rAR2X/VuhDbjZPK7IvuYiMtp9Nck7DDUWDkEmdX20ChMViW/zuTqDKqX22KFKsWqWZkhO
tq5vDsJOK/vkRvYo76IAJ9Wixf9lvPODVKPRXXqJ+1K4744J3TcyIOW6jHTMKXk6nuNRoCHWyxgV
+8nFzRUsxGQP/A8A5HHDbmH3S16JioqYxS7v/3jqBFe3KZlaoPxfLCoIFXsN6jBoQ1tKNm471FZE
lUKJod8EgDj/CMXfdvlWminmsyV2g/d4wu7c8okx28VG3sj/t9MWhDZ0cFmWb4tZ02H7uGf5k/9O
2CHHYqq3RXi2XJC1Qx7kYAyECGsW7IIlB3F5lkvCH8GaxlaoNO1LhdFnbnRCeAupBj7MLUh557G2
T6Tl1ivBwR/gSqmTRYtyYS6n7oLsA3DmqrFaeZqflFoYIXKWRJp+HCN7oF9Ktgd5+U3YDXs4wzLA
hVEW+mVoZZcvkUXUDnO3d/FA/zuXpcaavCgY1DZw4c3ce84Qk/gDgNikLUopgNOzkfESFrAPeOdP
8C4IOrHMuPRtqfANfjM6CrLeaNbT6D/Ih09kJcj+mf8VYb9X5wG7MN1PymFLT2BmAACo80U/MUml
rl9obhnGCfK0pmDYj+s5NeEvxlXma/FPay0OmRncBd+6TG1mkq+taXBLGuBjAxfhYtNwx36pKHD5
3zKYDTAV8C9dnseM9drGncDB4f+rwGoq+9DTmJORy+k4aKjCUM1ifM//zroB2aLbsTahs2Pn3nYQ
TzYA6ORWLtEdBleUVMBhp71qxlpzR80PYDggnKNd8aRSsYHydZSYpqDDBvw+4wdQdZZYEouuLZSM
7ke+PEdeytxvOEL8rgKwQ1L+JeB2i6epeiAmCRmjVGK0tzeALGwpq4WdH8myz/VnKqysdXCJPE6e
/41WhE79dBo+kOs/Eo2AF+yVAmSREg3+2zGV/jZ2o0bhAb21aJeHvD2uLmG+6MV4Lob1GFqQaNE9
PeNMqaBARoDWYD4kPGAfy8uh+v4HJD9W87q9zmo+/wBDVMyIgIrs7Pj/qxRZU41i/hkAiUV7FpBn
+3OCBpxf6wIGje1dyr51XIrl2NxRXpAwOHc+MNeuLXXMFo/gy7BJ10UxJfjUsBhXZqy9v4ZP0+Km
pS1xde621B3Sk2d4aa88vGGb1axh8PLo0vkcwyDCMqkPQueJkisHeCZDOG0ovm2VlqZwVpzUo7Cl
F7KiHyg+u+Whx9sSU/ZurRSzUqHe+BUCWdtY/PUd9Uu9LPkAZWBinT9LO7We1M/xLL4syzlS/x3z
cakpGnyVD7Sc83lK88ij0TYT8MxBCeAso/7wNvOL2ISjjEJtQapipG964VGMFD7BtMA+zTsfQO92
AfcLcdVf2Qja1cZiNSVwh+zeWGwncQ/XzKMEfDYIq6WuvYJ2QucnJTdHkdtipz4blkHjWW3UA4AA
nC/paFvMbhpbPemM59UC1ld1RtROMdmfUCQAfy2zDAt7FKU59hNVYQ5Bj54JE+Wsp/qvP1Rk6HMp
WJ5JMJuXC81ljaB3SlwO+PwKmIPSXfCBFPPULqPrGGNmzJ5wx/sXq4+yYlOyCrolOf46oZTHbcO3
el3mGV3oTYvrO32UqLumoFgvY1ns4AXuQadVzQjLv2kvS6cgxyTjtUGXC7hpnaRjV4yRaX8nEyUT
7rUZyvuqSw9/k/9uH6J47GObWVnw+buIftRj4XImBiphE05e4V5RCfv6yu/akzrDWToVWCNfJqtS
0husG1zwpI7XZvqhCHf8NDnVfUWgHt1ewExRhGFTJ1fAe0dmTIa2il+ebWZ7IVyMT4hE8O358yZk
9jMCtGSXGpK+/v7HoAxFeWNZLLwzZa+SA1NRsTmcJJVT08yGVrHDoaxyn9vNk2D9cyNB5sDf2yUF
yg0cSx9EKBiykqnVvlZti0v0deF9rNLeIIUU5b+UL2Z9TqwrixwSBOtM10h0LeE/4PHPmevpEer8
UnCZO2dbm4qK0N36ilfUmBAA/g4H/Ya58WKhuplhk9bEgl307pb2VUx645KS3CHuyUFXoq4MwEVZ
5nRxQrE0gdX4q1U6J2WMNEkLHmNpqIQc/Fc1P9lYBhBkMgptA599DR5brT2gOCLYUgvMvwMvycwM
++VnHzNay5ig58jFujbkCiyefrNqIdn8G4lWWt1lBL4QX33taXPe8c2DnjLPB8oQ6+8BWUFhNZmM
ztMDFfa37ByKaUqA94mPz7EOhcPEhMx7nh2wtLWRyF0T7sFpp6SqLRzIdgt+T5zayyg4zBNFlXG5
vNbllyHc7kbLuHFYf5TAx8YIU7UQuvELQKmdcujb/xxpRTj4UvP+1/mG2RNUYA0mIz3CWZqPr71R
Qf0ttmciZ2IuBd95OgFwc5fTU9YYd28NlHV+WgJe+Sy8yJFWB+HkFwaU2SNy3Lfv62WLU7eCDkeD
eJOXdGvpF+Zj0y2AR6u2kirXED48wxgpV+TxsvY8uoWjX9RI3MyZDCj5RdU6spzaE9ycSnqu+vKy
ckmoA4n2kjN1GfAfPO+O7gSgOFIIxl3T5SwU/xz6df8X3plIjjMHRsqdLuBYTGKEmsYGcQEbAbM9
jGeq5x2Y5AOH3Y8jga0DX/yo09eTQChs2BlZWNUTtRqFzbecG39ebHJ0/0Ha6+eV1k5rMFMf3uQv
uCapCMuiH2uRUNSYGOgmfLbBI/Y8dk97Gnxwvpth+zhWHLNRbDOBPGxZUOnE9naD6Z06fdXIrha6
zxODCOgYVQFXwQ667i9LbJIv9ZSXwbc9sAfpGkEYjNCHLGmDjx9Cvl1xa82vLyF/g62Y9iONQ2u5
HylGp/tQ5+kVfedMgLfalheFstesF44aV6pCWRRzUDode/O6fVF7EIgNYcMH+HO3wQLw9Ex84hJc
JmVyAcoxzJbB38XlQTTK4Zbo3pEkGTfQEUrbASJzPL6rTrUAUrBBPubHJYi8IymQLJeV8ekIXYkA
Wenub9q+ej4xy1+ClEiSgz9rWv+XPjsIJwhefOjtstEhUwOcBwBwKL2dsu637Zv8pgVIsZPS3fUp
fe90XH16RVPY8YDHA0ENm506byhlFNQY6ZgmR+VsXmLZKGQ8pp1Bva/bQ9qp21V1CcVvFX35dUa4
yKB4gBK6tZoj5G4PAh7ech6/APptIOxyMvP/A/rPv7wOn6DLKNZyTZVahGIT/t0V+z/FFsufjQhs
wqTNoFiKTsgG5zt8S74R5j7zzlk6QB1rJIXFsPBA5XuswJJR1gi7/TTMNeX55w+tkXs0qUO/aqcj
GsV3gfRbP6tgv34+L9dJWAGYpLFJZfYjyw8qTr1BkiP5GzWt4KKraOJYRCPjFLlVwcGPmJ4uBfq8
BJ1bKueJ3zJc/jRuzVx0UtmbdXCElRGyX5836t8fKXRXi4qeX56f7FUopNBadrjMlwRpBv/ACZUj
c7KIfDu44QoMa2DQxmu0tPbE+A6tl6/IksK77S54ZhFnrA7IzjgxTLAaU/0Frmt0g68uzh8dJA6K
ZFlmHuWNCV27f/wxrOTBg8S8nS1+jiQV/5gxqNXh3fKZdv+iyoh5zgsAqboW0EtNLZAJBOs3EAyu
z6MkcdRYpgoJt8lf0zRAZq6JtZv5OtEp5RCliqu4bGcIzuSp1/FIDyrB39VfPjk2gAxYpSK342o+
CqUOdI9YEPAQSUrtDAgMnHzB5APRlD95iDLxO4GGsA1nXyN3v0ijxy85pS+H/LXXjdIT6WVByl9T
vV7/IK5K6YsQYHsqefIwOOycFjcTvlfBYFh5Tt/1bdGP+oKpcYJcMK6C5Hg8CBckBe46KFVS2S82
kw0DDwfNzm7mvg35dBZTSjUOrM0dWVGE5sq9ahSvTrDlZ+9D/sZ1XKDx5dQuK+NNr/XlgDdJ1lbB
q2kutRmrXoZcV4Xxw95sBmK6kjBfWxj/TYNFTkGPTe096ct2+VuKr71v3KcIw8mtPF2+YghcQ0CT
951e2xn2acAweVejWpj19VEb8hMVsNWYdcTfl/BiHhxo5IpgVOy9zKgRzdWFBj448+cjer5OQK5w
l2iIzTAUGq/CQ8evpqm9vZtcb2TLkNo3R6TelaIOq6CXgpNGUZM27K1yqcxeqBOEoBh8Q5ynJSAf
pkGCiYcLwohPbMvpyAvi+HfMFJgxjzHLSvQCGdWwkPZUr2ElWe1iiodubhr/mRkgZR/gsEyZuUJt
9PaZGRWL9cDDt4Iblv/wTJRhDkgPu/GMgmhaMNh5A3FgKu1ioNFJEKcHg86ghK/tCcV/GPMiqPES
rhhYgR5ACGBp+JsyQ+gxg5JuzylcGZi4554N0uxUO/zeA6dKdXIeN974hEOsnGabLnmnL6Eut/8s
3ZI0Lvmfqx4r1yPAZld74wV9kn8GT7WwDm0ZD4R3yYBLUMO5xpPRoMP3kBGL9PCfnqPDjrIkvmlc
hwZ9O8gISmVipxwslXo7NVHJaRLzOuBJBKLpUvfV7cQGSN40eO9eRiOBXGFZWahUJ5ApNacKZdC2
CrkocliSXxvuD7/WQakXLuPLXayQNb9+uFlYo/+MUz/Qt1iC/LeOOwddyTaEwBlZd6+/KoPCXwOK
cp3alZZpLNB5qWrRgVPPB6np1ECcv79RXOB1DG6YujUSAmhGKD7HXrfPFcFGdoH4RIybtOpQ/Xw1
RfeO6AzKypRIKIdJHWP/MNKmrjqPL+QRDeK+xNXVv3Ko4UCiRqK7ye/E6qRvvMsYNvW98vEjw/mX
PVfXkF/0/ICX5db/WhDI13iffNlvw66ICQNXX37cvFO1EX1ys47pY74ioZw0AwSHjzeTlQHWVutI
RaPO+seSEgytRocKBZ9Ha/TcW18jQBY2WbliM6XN78greNsYXRxIPQurfXDu3mb9XfX4RnK8JzeC
6EF/IIMT4kjk6Cam3auhgh0cx4Ka3VwbL8IGwYwLxpUcjiiDU8xpx3nUSULg+f1//Hhs3F6E1gSE
Hzevr5L1MSmgYVVwKSQI2OGLc/6mY/TgHPj5LtHzOzaoGmAzWsyw9mSUluE2hlPqUdkBaICiAWvl
3C/Qw4jJsuaBFiYO0hCddD4RhuBuRk+TCZ0Ep93THDD/XxDvGYLtCbPxXpNCaFOI4KkR7ZMoaNOv
Fkp41/2qwpRXoAg8PM/g+i3Y8QZMS7VoxXQj1RAk18WX45mu8hZySc5+WnRv8gdlJz0mkB0dKCls
OMA+6kazBQuzZnAntY4TMt4hazEBYQK0/L6/TEP8ufQiVFwZ/Z14kojbalWqVtfsV9KEiqYjtEv2
8qePSOo9pPk5wZ7UW8pZFXLWUeV5peh93FHTM17V4LJDcvcVoGYa6KgRxZ+7DpBwv+SwO4dw49mD
W/+uL0Hp0TRJkq2kmfCtmVH2vWQLmxxjzA6MELh1m8AJqXJ2Nygg2pWcCHt56jtfZ3/H6qA+QMed
bHeHPIjK8K9QhnCcEWt5KY0cm2ibn74vSOQO/qehoQ8qI9uGqGkneUcQKkl7IQuYQjWD/Zd6NkaX
29lLlYBn8/2+fVIzzo80ClZZC7CzDJWjJLXFt5mlzbojSLNUnWsY7iXsL17QUDQTYg/Uug4TdeGf
rcVyZ/3b/2lJFcD4lI3glBPQ9K0mIvYOLYMlAmKz2HT4rbWNzXHC3E6WjyP2AedFV1OG6g6g5XwL
zf95NR/55rSyii83oLH26/gKtW7v47ip1hhWxQ+LYtFsXtiuqD+sbOY3GzkSxgSKGPMnWtNkhfwe
CaXvqkFdbmQvEGy0RZkQWLKV8s4gXXJhgcvqpm5gCZblSOj5IYrbCADhue7DGS1zfmri0SibutMv
rrlRo9FpyzikYciLWJRLttw7COP9xqPq//Kt5ONNCojG4dwWzllB7C4sHdkSptx0jRKcJ4nM9f1H
SPKkgE14h917CYk7NMq49ECmcpx7VpOrgB6gT5WW2XtTuMyONA3xyfm7qbwMRqZRrHtSu8Twp6kH
W27VB43+ZWBBi86PaVh1tZte6Xa2M6xzOSJ79nNqb+zlcoMGfseNE6W+Cf8UnAjnotS+zc522nFa
jGa9G9ghxzh19ZvBNkSHpDtc0sGDClMVqLW5kfaZVGLE2/4FB5kh1aPL5pg9UA3ugbpOar4YvQrG
IBWGj2E9uHXfPkzdftpwuOEAGV5RJnwJ9n3UZFUH9KRasuM2BR61pyD1sLP66einnZYno0RRPqNt
Em8ymVDYYLJR3cGF35bNnz85WzOoQsTt5NMH+buayzOMxEnRYhGUgSDB1aydAZf/+GH3OjGka7Xg
Ywqdk2ljthm2/YFy0ZcWw9DQewH6wb2W0yMYDA75L8mKAaelyMfCPd7bDBqbG7ierj576W77blr4
xsOZVsGAeefOAdSrxP8T8ErdOhf3AQNlhE/iHEWcNSFFBLei0Cwf92c7uTbUpEFUUcp0dER+A9kQ
QFWbA4c8us4bfdFcSvF/yh4bPMA90qZP2OZ4lPLouVN0yZxC5DyF/dziHetOvnDb4nnx1r4ImVPm
4TTGecFsGA6HjuiH+sqQA+mAeu7QiUA0sK1YS/jDC4EjCl8sd2uWLyohJLjWhOYwk+KpYUpWQA9y
n4tp1B+qVcedkfs/oKyPnQsmE36fjjubS2nNwW56fk3B3EdIloTpCn0b2gfXcNu0su9z0ZxQz2KS
prYHOdPT0Qnze6PxzbvA8JPXQbCdS8rKRJn0dbhHL95OkmMB7zGAy1y7cPiI+hXR3cp3ko9eHCDO
lBKQF//tHdZYnvAuIMt+Y/VPGqy8+mSQLWhk3LviB9LriW2Y5Ffmf1HnOsqzU73RqDDUec+2WfDj
nqGWPz5NMKpEYypCEHJQs5TM3EkrdbQoDhGWYr4yLejCvdEv0UcJE7R3eisjHKDLBZ57m3yaeHU7
OnRzKS+C8S1/GcbIZPMN0v7a7MRCxm+IFdfnIjq+PIXnpFX4DEWLA2KvySGShoZ8lw0jVY7opujH
4U87IKQym91CvOCKZ75CyMgBw8KJfeFLmvpFT3MFDoFj/cSSn3OnDK0f0iB/g3rNfzpPOEu6YZz/
OTZWkWZZ9WPLcv4vFfx7R+metrGMfASbPEiqSwBCJhXnuxujsvoKmEZ5B8BAgbvv/8WyppAmlYMm
mwXakegz8p7UMNTVvcK3QD81gKrBW5/IHYkXmUSDea/OMBSxV5v+mwWI7q/7qmKex7bREruCLDd/
DbkaH40YxSoSmErpxowksUpcF/KqIwT0hDi8E8vxIzR4mLLGD8c3IsV/ElyUmDpJMn0ivgIimp1O
WMQ4PfRVIfjOPop+6zz74bQvV22kgGxfUW1dsO0LwSd7ZIAeMdS+8bzDTrKGtTjlN4fqhxePNiyl
cylBauGdnu1m5k3yPKsf8kGrT93GSga8cynbkcLFMVCQM1TBZhT1ZSR9ztw81qMo1KJBfoYu+NJl
uGwSeba3DAtAWcBM8cYwz4GOTbLEG8VRMfAp4iZ8E2+KUJao17H8kW6RkuMXDzxUwE0I1Uu/KQ7C
6ASLB/DgSMC3lTftP1IFWOs9qi7KvJNWqLS7SDqyt6Sx3PLP8x2LJbhCJ8EyjOgzwBvHs1tpHHwl
/x0uneIoH3CveaPhCcmXNCCuiCYm+XkDBGBDJjo1eWknw2IXAFyNBW2PPwn7lefoptkipDefIBYk
6hWnSYeKN1TnlZqMVajNmrawsHJlIoyPROMLDYipNB3KramuqTIjySx6q2yuHITfPr1H2Z3sm4+6
IyDfZgnCe9nIcqj3s/kdEI52eWDElsqE0WuyC0MPDMxpLvgBeUhPe86lTYMtjllNrxjlADwpuaIS
4Ycts37NIEM1OTGlKtvJv9ign8wG1QiXSIXec+YKEPngpv9PJU4T/bsH7kIvfL+m6RJuVwy5QFrg
QFt6RiHQ809LcJzY1xY9lEQtAKaWx4XqXJsns+QpDzgUonxL4e6MKun2VvpSrhNe1UeawjvjgdiI
xb/VuNGhCp71/begyRAbzmSRycHvDqH9riXMLVp7sSmLMto/4w2aGei0lqA4nJRMToeNo1HyPTk+
8EjpkFI2XtGV7yP8NQr2Z7L542PJFTbjLGDcgFL1SvwDe/XvA7Uo4aKjcYGe1LU1IW9fAn+QM7JT
B9hittDZUtlEcag/u3J1N6VDujiUsxzZ4ClxGOLZx9GVd+V+Ar3x1YkK8/plbGqVmWtiMkJ6mGD/
oXHl7Na+QCMSP/p02dthehQaooXfQZv1nAyU6xzEkYaQG52Dj6pDk6bh7XZNLImMMTI28Z96MBPz
gH7jH11DLsEmxPMutNFeS1iKu+dUvrGh61r3GN40ddPemUqzE7EH60vc5yZnj5rTs9h2ZzAsCKrf
4+2hiwWuLeMdQSpRDBIg1pIQJszaJV2Io+jpNkX0/Rv431AkHJWMrLIF6Ly+QOFYa+hJSVzKYquH
QVB17PuLY6WDvzub/zR4nvAhwHRq9R3cTHQOGp3YL1y5N6iKRm1jSD0RWWlQieOlfSbyGxIoMdsK
9ytMkrCkkIpkSEBguJvIorXctll7iZ44WXN0VVozFtLGHKMvEbLAyuaHe8IaKdvUscmBq2Rac2SU
vlC5K42kGWqkgEIHDQVvZCyaX0FFoFCLHqa82uAGQ/qs1ayvuFES7VJqmVGMSbTQKPG7Bd51omlr
eiJtGyiZBA88V3aNagT/++2QAWEUhIdifJwMJidQAjzrRlfjdoS5dH+AvueDTFHj8qChwFBgc7yg
OSGN65CJPBpoeCCvQ53xlE0x3yWT3EJWvj1e1I/rPD879EWvJnjACL/paKIxfj6FPQj9M9vJgEP+
BmDdZ7djxptHVJ26TtssuI9kA7/u2JpXH9Gus5IPShNQ3TesPrzfNG9DQIXPa4Qg4KVZIZF16oOl
oOTwBvJAH0tWPvt3dWdOM0HXSQ22INOZvncGkGmdcSFqPPL02zdLgZMGQnJTHPh+4/776YgF7frV
3ZKIq5aXCnmWc7lSNPMU/6xO1zPjM7JwJJgPODg7r52jwsRunjLZ0qcBOKzOR3CAd6vZfQ4IA1L1
RGPUFYbiJkMtnVHpe3mMffFHf3o3Dknt766b/rdwEMSwonEiF9v9wNdIAHVCg+k0OLbSG1MuS0vk
Toj/gkWWZh3dBAlUddyQ6RbGlDCPeKliG9CO0i2YxZfwRa84pcWbHXTc1BB8+3/bXqHAt2ny/b4H
NJ/BAWeQGWjALUtx0HdheIw8sxm6Opz5De0ZNcJyUb7falzR+1QeeE3eVXkpR9moOf6sV8OvLC29
7o1cAs7GZgih87arEeqmOJfrwqsTb2ZOufDARKlARHAOUTqJwW59tXMX9qe4c1DueH2JP8C7qJEs
Pz+G04HbeQRWr7TVRZ4kMS/NTtDnXEhJaXqqNcJN8/rCEhsVub6ShP80mvBu4RzoWmzlQVH3Et6G
GEwl670gvHEvHuLPPKp77rAGv6sa4mQ8oQdqWWqBbXgSLUlk4nN4kWdfp62e65ZbWICuXtqxauiW
C5oADA22acLJmw2BiDMp6t53WJKiXsIlJzrCIFaqS8tMnEREZBNp9JhH2Wztz8XyXbA0nPr1pFjw
P9Hc60zwrkFMycrr7nKXkjHzL2Lu7OH7TwxH8rSoeqvZa+O4rOd5Vn6LjHbonpovj5wqYizfPAri
TIOKbxAmwczaKcSWGR6ZOCInZNAD88Ago4RmxANlkFT4Kwy9Vds288OrwR11MpzRiiRQnntlISBz
OueleK0GvDOQ78Eu959nxfMJkcmTmc7U20+A1IioIgRgogjZ//uRuHQA2RLRqL/jxBRT/m6IwJd9
CRb+Pxm3N25L6FbVit4p1eqkso8Bfxm1f+KQpVgwqeU5GfFT91L2kFW4lZLRT0ck+oOy42hxDZdx
YabG/DATop2kNq5XdSuBgRijUZ5I+GyAam0LO3wVGlq8PPdOmD+h8qSTUQSZAf+wArCHCKZGfdQf
pxLvZD9llJ3/+gOMXXjQVN1pHx8OZUckBRow6E4QVdy6+eu2rYwW24ER39hBiACUDnMNAhfHyTVX
cwJZtFAApmgOTJ+vNUGZjIeRy4v0toAHf4HxtsvRAdJKfAu2hnOSdkX3IEXcGqovTCBtVuf6BzL+
se/63frZTOTryYnE++80nYSlGsEo9zGns2+07imPForbEaOkEQYhPpO6RD4jvKCRfuera8W9jiz8
nFF6VKD4tm/W7esrAy0oMiLPTiiI3WhHM3odswZDBeKiavpgJRjkm26mrTri0WOo5/nBI0v8PUVH
lnVOumSjza45XUd3FPq2Ssao+luT8gaoy2vGV7vA2OjF0YVTtAnB3RyOSvZrt3+T7FX0UtlTxvn0
2JXLpkc7LzLLF4miIjq0pGBiAg9i7kE35cztCg2Njvoi/gZ8rXJnq2H4y/Nosmg8EpmP4NfHzYT1
9Ls1gEb/S+k0sgxsBfoEa0MDIsRjte9/8/+umo5L/1apvpgvDIJZUiutrnyDfSdQUffBsldUmy1i
T1nFiypAlCo0RX2wBgsEnIjCAZn4bRHKjre3a5LHXdHLRouGu4eVhH9vIpFkb+JcIWu4718gEac7
NS3goxs9/tG4WroeM3l+DBMJws2hpVN1YVo6ap8hHFSiLbiwuTkJwns1NEOGTqgq0FIiiguPArFD
s2dDS1Cqqqk4m2DDIA2f2jBUJ31xoYNR3IcuSLNMCGLwlK3SPxyq5ne+5D/vEgNyhuyI4V4Xgapx
DhbayAgDdo9o6M9+7dMVN6+63J97oDMv8U0BKp9l/ekVRD2CJ4fSSfLThVpAncgUBkxa3VFV+xu8
hWTx5KFe97oJqEyyW8Q2+QV4sJ/yuxzOyjiMZnjQJpnrQYSK3XosxyqKZubg2UN/zr73mmbW0P60
0CGUUpA5hmHa/39Kl53o7+5hSEBDg6/SVzl2DS+pzNjfhJ0VXxD1wLBMVWOfQ+1F1nvl7NoNHeLo
Y8+Qd6bPajVaNn4ov1ePh1ubBdDETCom2d1MIpDS5w7nfWoZ7aOH3KtuirR0sfPfvxU4dcPu/CMx
Q2rSqYTomW8ovN7Zdc9fB2uzoDe2+Uet7YKANNS1nHG5+s2uo5sZSXKzCSeXUSY6SuR7Gsmh3yVu
J5+NjDVLiY81rQjWPYfDAk7ojd/LMQMk3rq7GATrD7nHGX4fpHUWpJRIYDrtm4vXiHH/M8AzzqnH
4id2WjtMY2RKv7jgNHYYM6H8V8lkodSK/T3IICzpBWRnNNv1BAN55Ccabp60sC8A6cTzPrdXd5wW
kJBgUpb0kcJqVmiZdHBJVJFtbmzGCO8WJRm0IMlAiyJR58dYYU7M7WkArMr6dsKsL2dhyGGRPPt7
ub9fNkH9gseiP414Jdqh+1LhsZ4PVK7pmTCQW6TrfuqwGWFUE5TlRDneczsmNH7eX61iMsZNxdbt
hhUyyDVPJzx+OzZ8aOCkytuwv68c5/PMET1yEHGD5oSEUHTpEiWrhiQzk5UF6tTFp4InxTPAWfEv
LG1QrnxnEYdSLH6bRyH1N25J7sQkE+oaEsCbRbkX7SuZErA1S2CMOaVwPS3I3pn5QeqMdCRWMvp7
z3r/j3UcgLRchbF0m1FtapE85Nb9nCkHTSZCvN4kxLmMo+KiA4JSOEDeiAj8f/XKKHCwgr0ysLjj
OsBRM+DPr6TgCdFj94PzzPa7Mj11jt8ROp4SFQGyRVcn72ZheUFg51xovXaev8lA4hQfuWJGCzJp
0mucK9nc93zKBr1JbRSnTZhqBlFDqvCAyllNJPgkk9scNwuNYlMrh9H6KVYKEbwBB7LyGvKmIWN7
4gyp2azvbOBaT0siKlAm4G88iRXf/Nb7B9iecDzh5MYBA5+obH3AvKgJnLeYknRjOjtwl09Yx067
4eDhmS/J4JcE9nNLOeLQ1Ao2ayHC1J/yaFmzSDRw4boTXp4/fTbf8vxzTR62tX377FhYzDC+r7om
ELJ9Mr95acqQuD6xK87kr01QFBdIPrpuXkFBkqHebeBz8d5A3GLldmLPldNiUqR3Tnn99lZ405Lv
e9rhLH9g5lmOocRXhrFbwVO/LNpztw+pL9hCo8KI9NW6vgxViakrjlwxq76At9CQeDv2aoS45Gbc
fOvSfuuSKHpamGX0bSgV2kayf5/JmrnIA+NWQNE/SpLQzvNa6xPioUjPvO7B7hoMUlguIevgW0kP
TDo8+SqLkhs/NxrQKV+5dmjX3HH8sayYIQDtAxncz1XovR2qdMA1twcMz1RP7HOBWq0AzG+WkJcc
xU3hu6Nylo1l/GgsptGApvtRLjT3I0b275ggfn68igS2EfXkIzGORQP5fsxKOcCLyqEj/wai6y7k
tGB43Jk9ia5Vy2T2dLulMVJMpSqrYwx+qRYbpBoyDqwSxb9tASwhxtOEQZ57iBJwWbbn6dXY4c0H
NhWqnr0IMfXpWq+GeHQ0uuOiDtw8jRH1itK1c9zPW3jdEJZa39X4QLLn3jmL/D3oDK1+xfiKA6Nn
hbbJEcnI936BrU3Pt6ap/B/qxjm4psK5jv5Bx5jeNNY0VWAwWnelldFdqgrWcubC3xmMI+wRjlh4
1GFKqDKXfWn+0yL98N/RbHLZV5EV1sFwmgcnT3mbueTdRnE2hJBXUNxNRnrUHSwda+PfW+Y8I24z
4ZyU9tghks4+cetuzkc56QQS+PsJx4fVZXRsKaJ8K6DTGqWpxtM+jk6I0oiNiHaNZfCXMVC66K28
6ECdn6mrLs09bmELBPT3NfanaxlqMmIglDTziFZrehtyhs2qw9/aylrfKZ1RpZlMNAPZBIyPM+8a
isjSeA/yaAg1mjau1vxNYa6a2aYyaBphCAPSmk2rkW9UCRUa6nD2XDt7QZAKfE0MHfJVZZXp05/d
RW2vI02+uDfzOz6f2EDnxWXhFa9uTQh1Tm2QtRZZj793T/XHwClikpkIEhqpxj0xzJKCfDRP2N3m
7RrEJWFWobaIr1wUnB8sT5KBeVR/ozcmBVh+u0Vglpy8lVryqHY5qAgQx+cAeWTMXB4SkiJlnLlA
6UzapcvtMbxdWlC0YlWUn+naecHnves3jfxiyzdYf/Hbmwl2DcDh01oPvSVW1wnmgdmeu0iPHI2e
cuIghOvRhCzg6JUZY53TR7yhSWgwTj+TF34ouHGw/kXvHhiQYE0wKDaKtQXlk7JxvSxbqLVZ19W+
605Bgifdo0UwA7+tGUlwkQ88qodDtB/7Si5fZ2ZeQwfFNF/wWmzIJA+yjar6123m0NG5tedFbI/c
YjtRvZUwmooD+L2tlJlowq/m/9/GZnSFznjqd7zeETHZdqzmGxK4qdggXfxccN/WEGXk5SYZpJIe
SD7uerK0cr1U3Tffbgb4GzMVdqsKln+Jj4mXOCUMoZSTvGuDBgIx1fvFoUdhC9S19/gMqMrf1IEG
hbXGHS5rR4eNcgbNykrdc6z7GUHMd1S5g0W9m/wUYsaoYHx4xR+86r1EygCfg1qcc4bM6JVAHyrH
U+BrKfWQHiyznft2G47F56+U4p5OAcyYNwWhOY6al8gxHbiZ7WexQolv58HLnQxGTYDGI3y0HL4A
3WYdFzX4yBc99yXqtxk10EaCjxKEU/dOf1e8APa2ZSFeWftz5k7wA94mH3ukmYF1CUOFNRS5Q3m5
/aTuT0Vn+TOTs7IFtPX+DBuIz8JfLyGZMCD/9xbLJY2GBHpmC+pOrXIkEN5afVRv2/WceB4VqWBw
hqZfsohO8XmVL0rB/f7jSK8QLxwmJkRznx6pW4ePHF/pCyZWdQYzeQQEtIF0wFE3Qflx/dLmrTd2
A1YDvf208zqBLcn4lXFgz/hkGZloxmyjXqdPUHKZpLbwwCeMtVTsznmJFd5BA3EEz/AiVNF2MCLa
xS9hrUhOVgrDhmW5mDOvoCJb+f66QgHPJH1qsMSU/drQ8UAYf4AaiFQ3jedpU8tHAajYqxg6ImnZ
J3i9xtRy4q4dOstuB60v2dN5oNr2EdYjSoSZXRaqyYTIm7MxoIdP7szV2a3ty+dg1jC/DvouPnuH
dMezw29GsqaRYDrGcbx/Sz4HvAJy3BuVdCIcb/QZbCG4KfoR4fVFgFjMDH4p/NIxongzLKRaao/Z
2vc/QXV1K98bwwGJum2Qd8U1FAETWmueFmXw832B7xqTadBcFbOfGuIzu9UMr0sD6LgvoueRMmXu
l6wttSbfPs9dssYj9WQA/j9wVdYeQuN0+wTNqIbkft5duPhZu17TEHs5IAjgYC0oWJ8GqyfcfYP9
8Mo/Mr81SMc0jsI5SUpZ+KQYA3XkxMuFVSVWeJhdpeqn5NF1Gm5J4iQ+kAThFwEY2CqOUqEmSwbP
FpbJmLCxEwtJdbyQwPtm4B3rS/u3Jr60liN6Jh7ZQsIELkjHWXf7Jl7Uw314MZNc9wtYhVFzcN5B
+i0j3GE2X1lS4vU8o3kecwHOdPylMstgj1/yWfAbHwBvsjgW2gPoPGsxRrv0XEEB+P+yYqZzVBYD
X8GKtN4axpXIZpmTIeV/5Wp3RNChSMWTYdqK9tDw/GW9hqOKk5Az8Z9AFOZeRKNLEDdN6aeoLnW0
oDE+V85V/Er0fDux2mK5ovoX0smjQg/Dykob6z5hcrHAarApg8i04sf/81eQes+W6UZRcR107bG5
YAhVAn6OKkZiDcqu6qcvrlbg3IRgL0B+KKdkcwxPWzbFzbeu+Ydzr0iEPkSpo2U7V4MWJ+vEv7te
GGV0n8qKPryaJtOu81qoWRqyjcirS/4O2VPnaW4lXrBHlPLyXo1PNIgBE0+3p8Spxh4rwpr9MN5Q
Lc09454qErku+NetlzZX5QtsqRIOjVGg7JKlM+NyEgCWZUmX5IKXMu2QdAEfxb+PDs1GzAU9j07P
uoCoSJg/gyBrBp2RlcX/EPNwneie3gMBdEUrF3duqIBHbZ4ABU/aRtlr80qAShZhp//PFBIR2uZr
sA+27lzaJb6aviEYPrvVVCUSKovSBPfs4N0kDXU7XczjR5o+x9+kWwmOzFpGVh2nMCw5U+y4qHxf
rcfr1kMVDK7JBK1ZExvpGEQkAdn/8DgGUcdbbOpL9rx7SPAuQbckfVkYY9705kRl8NBX2EbEL8b2
gwm/rJj1Qf8zTK1oh9yTTYO/oLvuK23xRSlfLeJg5qnCfEN/ZnKa+ay5XT3M9p9tpu41PBrRf6G9
/EtT/KGhqpNuxzZxqKg9JzXV1SmwaCFuLoZFliG2gppBeHWLJr+M38TYLk+GzjkhE0odaMwOAHOf
QBXKgueA1IL8BE4v13w9KjOVblNLy1+JfT4lmMEwJqbpqNz3lXIUHzkv3mAj/huP/5u6KGdXCrEH
mVFOZozaLtuFdnFfU0OAgPa438a6y/PwN30/6DVNFMcnjgNqXOz8l8/Q9J7g+WqFFG59T+AW6DRd
5CowIlGQAPB8T3zYcmwtsYCLL8F1r16POFLVYch49S5Z8NPnclAeZ7VxoGDe2nhKNbMY3bYfM2E5
TtXa/YbWWr0Foe2cmJ9Tf+taAkU5T9L0K47daSjF1D8z1rl4DruxbHKqW9TTN36D4ZsLUw6nOTED
QVXSrMqnTrEGywSZnDDAZq4awwPrW+Sn1egAXY/pCoULgMVc1O8cEz1r06muwY+Pq7LgZioBjQae
TZQEb14h5BvY+lHqxto7frheHMoQqLfb2MwRSKf8u6EX2U33ExgwU5MkeI1++Gi2ZKdL9ZB0Wb2d
LQde+n1tfNWqaHhvdpAbdB99bfnPZo6TsGTot/AVpU2WlDJGtwJy/43xJAWfW6rRyyPZ3r4HGda9
n+FC2H1xlBd1UM54eUOIDaQgtIadFHHRzp6yFgpuJQTECsHML7739Gbui+0cUuYKQRtHpmZ0GJJ5
XOt8P8f5kbhLAM7n1lVBsIFl0dOGw3ARBxXNKyiaWzJ03x7Sv5CdU0K0paS0OuJXVxfh10quQz0d
+sdaFOkMsWkdPe2BnYEvmFJt7D4Xe6QoWRlb+gs3F4v8EmCnlpZdq96SO0WeIDCaU7JYHPddRHB2
6eX9AFTzY9in+bZylig0c3dCyTxIfAWajv+AWS2MbtwL27qEp5efKDujsx+9Th2ydRBMPDYKi47J
P1Fm3Z5Tf9Ub6GyZglNa8GBnZnsxL8O51oasWicD6gL/Ia/esrgVCd2EDr9xCP8MBH2veap4cTXw
tyj3X1+jOI8ea47JcZRHuNmew1ohYERGXAbEGPYhFnfAtE8lg0mz/sNuys6IRubHq5wVtoZn7eg/
mL/hfq5o+IEripGsoEn+z4ohHfA4CWwEVxtZPSFHAbBBMr9cNcKWhhXAggsVYZgqEUyxaefQT+VU
OMoLiUvxtQXv0nYIIYv04kmPlL7NXvn6JrPXAmJcCitaFL5qhB6ar/5MQrLhwfnnHOTqzFJcTVm9
cZpeIhNIF5gP1+EZzrYb0wpTUh+bV1+yy8nZMuOVOFQXCXQpTjLRBdNsgI9pSCmRdUW+M0OBvP9H
k1sFOas1CXSfEgPdyr+J4mbgx0+VybcGqJ6R1tBISU6NJvzERxN4txebvFkeabII49DEfEuzdr2X
GZK5sPIQvGZm2JZM5AXi1+FJ9jSWTlDkGlmXc5foKbqiX87PmEd2YVUp9QwU6/2keKqTkDnlroht
KY8fckobc+S8rk+01izPwuIpy+IFy/roUkN4KVz5EwDmiRI4nzgTmv6urIWZOQbY8viDZp055LLr
RdFFEnNBPJViOqGOdCQj3rXISZ7IQodd/om0x45x1wx18GmInvlci8VhDyoccqEsjfrWmIsKH4Zq
5y6DhYUkaymAXQbI1BPQZtAlMjEA4XN4oLOFfAUvjncss0KRFGwUno71M47ylB0bAxx0uMB7GD92
tE+IPZj8T77L4SAUnF76e4SQTDHITMO1rMVCJVua9e5u+Kq+bZCl0f2lwep8QjaCiRmxe/DAGzQn
WCSqg2dfD36t2uAIq30aTggvS+5fYeuKMaRwO3pLSLc2tmPqsDWwGdQy/1KCkC+9scNHr48W7BhB
tT54GcC5x0qrtfQT3gX4VDh1BcwWLApDZFISRb+lOOPXu0opBGKBAY7rjolzbxXF7k4zPGBlvhUF
irmPVrM1ErUvufJDhPVsZKSeRpZRmjra4ZMvzRsxhNXjJMMOo7XaQMsyMncsZus95xQA51SMeZ0f
nGImj7WMCQXdY3I6FlNrCGLdH+Ase6cEgMLmV7lRg1Bb1Iuxx+VoTE+1jYbMU5dmFHE+YQ/8/2St
knqsu6w/p4sZJs0wbsumChg6aRlgToLGTwUPgFyB1bvfozQcTOlenyVjFib5BUbDfFyiDNrVv7RD
bws3I7pFtxjgu4nX/zPYt4KW+vZwdw2I8D2zMDd5R2fAfoOEeVC7LwJjIH33/CiZPhJVUon/wLFt
X08wtUQgvkudrxNBFXmK6LH2STkMobwyCGGJoqDAIdXHeUVgkAtYlDOSnVCD5OKr1yR689leR+JR
DAdFXV2AzYeq1I22hC7VN6YPV39xItrZpHis3RuC6YU6Gc6stGRkq1+ElAY9rJ0FJgveClsd4LVy
cykXdx1n1mOVy4+P1MXIRlli5aewxY19xjT1Kj895GHtgMfD8pfiytzFkigJzA1+RI6mWa3KSaPW
6iwTkf8X3yc1sN4Jyl2WcmmHaZGdO2463GzPf0OgJYkFL91nt12d0TqWErF/jkBvm6e7Sj5VS1a0
0+ubOSQK8/0BTLIORqylgfc6VVFIAaPvi6gbesT+P3g2wAsKP9K2Wq8ebPyAfR1E1XT0cpyLdnG/
O2LR39Iir0bFUqz0YBGWke4uonO7+cvzsI4u6/Wf5EEd/H5KNcWBNsCUNRYj1pOod0EaVEheRdeq
IP5rklIm3ifaVNICjEbtw3Omewng+tkAvYTHgZ+qNNvdoyDbAOtm9/1jwmzXbv4pwIjVwAjapjGU
iDPljA8ioroaSCT2E48HtDWGAcYaIjfRi0d2g3S20Taaoq30zxyZxmfF7MGNrxfjl9t5nRip04Cv
63pyDnJYIgfHChRcO3dScM0p2KBiB3cfDg2car1sdjPSjHllOOMiycxNBISFinnX617CO1k/KNB+
WxmJfhG07d47ubtOqe3b3ghmGM6eznNFz79v72+fgfuotOO1po20tkD5Cs7NGNExEoBRqIVSafH4
d/BVlHozQ6Adj5t3FH0Qxit8zV8Aq6HSyeWm7Urs32+j1H+emD8FlTZVCqhoiImZcSblH5Yu6qGx
6HLnPMAi7uqOsP1roRWO3RwOHitNFzcvEti9nD3Ab7c9tb9BXk0czB84ayIWYEZ8s4lV5VLaH4ut
YIesso3Lu2lJycrPUMJ1beQmqaRobTOJojWMAlQbtuG0ay1v3xUmH/8xUCW9TF+Ez5zQvxBParAk
aZ7uWNKPcY5OGdQVDCoMeHGAWTPy71FIBGGQipLBa18/NiEcj7gxiu7nzwvYLsnNrFg9/WE1TwJw
MTha6ghyqkn7kU/tzQjEhGnl6cawfStOmBXNmbsKJ8Gkbf+4hvIF+PCiZYNStZCEgDh5g9ioNJem
90pQGuRikdO5vKMKdUTJ5YLL+aUk6H5BvSEGoeDnoFtTsp3DWvWaY9VD8CrvdWsKh0wZ1BtXseZ8
no9dpkYXQ93sWY5Y53uYQRmkYgs6KJSX0dBod/8FeCbRPZXuBFoCo2ILOsNqWP3cUP/Avs5AYo+j
Z+qRsZ9TM43Q83NsBp/wYjudqvDkBvs6umPuSN5/1UREf+IwG+X9QTifVMMzc7flRACShFvCSwUK
8V8AD1MS+37HI+9hz5a2rp3ZbzL0BT5OmGnrMOK1cEQKfidYQSuUdUVhlDidrbPYbFihfSk2n+uV
3wbgBZGB8d2g2f5vDlYxBY5g/H5Vx9Uhdx3iSeaw4sVCGffh33BXZaEeeAh76juaO7ENdgbIxMSN
Fxeiz6BbgnSVWJ7HFb7yGIoWmBwfXc6pzljBoXCqSU9YJx73AGBpqGALfBvJArkKxBP1fGGf1pJR
PNuLWlNlUxSU0jEFCSBAjhFYFhcBnNjHvC/0sADl/4UnGku0rv05IlnwykPDu5Uz2d2GVx/ntXHE
/fvKMUC4i3YHuU1HQWSjD6Wzg2MR6Gg5x9oKqA1YIyO6gLVRxshg3j1DdzVxNQECw2C9CVMekKtZ
zIXlce7HdT3f2C0oILRuAuiNI4n5TOCUQ2hyCB8xS2NyKYC9PsonX6pyrAGKZ+wSb5SAPgomr1Gw
1EMLbviGe/fQC/jr1IxWrxtXFQGGj5etoV8kml48iknBTqheplepo4egxt+xIIuMjGvOOGV4Wt3W
qUBMcuSjHa9xioiRsnwurmolhiBRt4qjjoQHNp953Y7InKYOOUbTRoO0sVyGRcC4wXYKDl8Q5Bni
6H2JN066bmoLYCqhskUJ/5QhZj26/Mxvp/R0SvFSm2289n6evjU2eClq/5uzcyqTVZ+bVqDY/3sx
0mFSitOCn9112Npk289leqwqyXqgzPA1Phau0T3nIJZdvXQSatv2ovRKqkEAUu6jA0gFxHQMCJrE
zO1rkjHwrK/p69IeHECNWbev37qRNbV+empCHt0Kg3C3Se591OjakJfPXZw3DzuYZc2Wng7Ef6cT
B1EP3Zq1wwHzbI4/tqJRJCiSG7lMZas8ls5jFmDg3XJcuClowXdg2STB3Kn8f2uZE2snlIFgqhdu
KkOmRTM1LohOBKw6jDsIWTF7iagncYq5luQUf98twvVCiZu4IxDnD0O4Kf3oraXZImW/90dvB8pY
1gGXlKSpdmUYcc6t+M3N/WW/Wiqxp0dWQlxfJhPjy4CR3RnC5xiWT8GobOCFl0UsVGHL/LfRt6GC
y7NIOiJiMNXTFP8huUrqYp34HHPsUub2lYKBFlag0N9d0tOMKOxUfUzhtmooVICCi/NKFR9i58RB
Z2Vv9aNq9/k3fmOhrfm/5002qNARU7G0+Ou4p02JmrMuhT5PjEV9VcsqYVSrTTJJXqWOqT5+8yQA
UFR6dN+G69Db/eAILSedIFkY7w/FaQ2TPlD9vXEJq4K3Uo5B1crrtM2x6r57L2yMYq6AJu9fd7ZF
36Jx/qLzpD340n+Vu4qo5LmtWoRjKh+pIMcbbPlZZzN5frD50KApzgb+seOo17jVAPPAsVRUuoJi
/o2LzxvWuq+oTciNBSEkqgNj2okDSzN/ocb3fhX9HDyE4GOctbVTsAHC9CgXS4jjXvc7wJJiENh8
VEqGqcIBZDNAhA79Fuk7hpqbPd+gKWyfoXQ8ODkb10NqEK9ZwmxxJaPNzNzaSVnWb/ULVgts1UYb
MFoJ8f1224VaSaCvETLwqKrTLx8EnuX0pHNhse5PVrMDE3zOLAIsaAJQbxGeSy19EjUPUhEPgbyB
+0DzEkEkq44y1+/T7kXyv6Rluz4lpUIaR/4lktab74Jrz41C37I1G4zCVepaxXJsF+oItB2dN131
sfzuBOp7DDZxzfyhgh+++9JS02+x6Rlhl1/PD2mjNyPpnPlmT8CfepGG+yPA692fgknBPYgRUiPd
OiWHiEuDzLOFmb22OOuKNPzT/K0xxZwMgJIvxmFZlV4q5q7N2JCrhTFyzWvNxdp9CzeunWtrovOo
O6m/cJvaq0IriyfT7iZQlrNn6qHe44OmMBjpkMoOQbFe1kBF0p6SMJDextxHU8rT0M6fI0NfODRT
DScBNGuFv++Kdt8eWJcfoDlHiuwGUsniAXzIY+4QTLanc2TZCNdVElOLeQyVZsg0NgvbcSfPm9I8
R/iu6TWALh015HyuC5EyizCHaLn0PMuD8thdXXpsbdLW5VGZz+/ou1p7hiMZ1sxG5qrI6ukQZgVp
SpKxjVATCloy5G82ZXB8rYyulqahFFH0GICGcuF0FkuyqxLzJKLYC+DqvAt5ftbEBjvU5mWsFVXN
lLtI001E9PYfjYQ675gCelnry1oPvkhs7UMLLjiB51lLUcx78hpFgxaDubHgk6ZtWRDz6M/EsnA/
/x2KQHLr09nl+w+UvwrN0xMuMYOzGTFnEdhaw413jlLClRehm9zphzo5UtXwR3oEAeTjbsn0eH9D
Q6Pj/2+mQUm/qcjrKqG4pMYXo/xrb7VFh7B8flRQ71Bh39isUsluXLWdNf8xkOjuGmVPxFxCoJY7
QZ7RhPjPE7ndkNKQZ/jCgjKgV/2soaKU0PGyXPHjPQ1tdKWL0fCci5hQDAZNUXlSnd6b3yP+69R5
azxqs5FPq+oZNWYXM53GxQfYR9e4VVgOyrq/zfZj5rWxpNLkX0GBJOap0F5K2JRhogHE8eXKOrWO
3pSgpU8rYrOJ9hMvJ3mLmVO19QVo0U6JtfBxap/sL0Wd0fy5fJ/JgHAABaGFuVcY+JD0JkA1o0L1
j0lo8hcT3TPcKJhVmhfoOyGxQqhbNUuwGb7H+uo2U6LQvZw/GaQVSWiJ9wYvazmtFrcihcXiWH2w
xEmLBc7Ez6U+w1O49715F18YY16ehMbVSi/QFsZIiMay0M6WE2zGE/wX9Jrt+Cg/PCcDvVbWLu7Z
tkef5NYDSVXLZ2n7Y9NXhI/eHYfVBcjfwp/5U2T63+7L70NAqdTwfJBwA3S28hL1l2Z0rwHJBdPu
gKq0wPWMuoIWyOlnW7Rf5MKu9u/GCP+ODJ6Qs1yHqtaa7lgvkxD38Zq+9jBKjnb5jvNfd0bQohSY
lEo9BnwWkecP64noNURVixhWpIM5wiMEeMztzmjdlo7qW3UndgcVFRIH8s/aMrfZH3u8AVd8xFwS
Z8aCz9K79y850Dl4+UGkLk0nXIigE6pZ1YkeTBVxPqk8hqvdpNfMbaeDob77VCd+lUqRou1f5CT1
khAg1LBElL70mWWrSUWygcAF0E+zWIV+nElCX6mx8JlOgMSmuaF+npmkRss/cSoJRzlujq2mWEzF
ay/n2aZ/hNNblUBsui3l5oIzYv4j7Q2t+B/OD+kboPLXTIRrBnxgdEgY48xCDcM62u2bV+BRzkjl
sHK59gEZnnRy0JHLYK0n86ZuWKUlblk0+ktoOdtH9KH3ZFjvcoB+zFkVwgjEpY8BxLN5tt/B47Jy
PpuGIA7Sv6jLT9Q4kGZ26SiiO33igjnArLjSqFNhEqAR66hzwJ129toE4W8tTAPO8mf9qjUgwfNG
2/dvP1POJeUrJ/yHWm00Ai8JceBma8MJytvQT27OGBAjAOErCly0qyJhsgmsFvoZzZyxlWDC8HkO
jqmziVYYPWFGXDUPQYWYHtFiS7tRABFriA7ZqijnoIDjdj1bTIp+S6jiKg+GsZ1kocvbfV3rRKY9
Q9rQlGOtyQSUHMpMGnJkljFjiKsljUU/EUYUVih0kNUWDI/T8MvzUIAbD8Nc9tqLvxGcPyGVcB28
1PeFktm0JFR0IS+7dCZytELveDtRrF9Q2Toi6V8e0yI9buIx6tFgXpa3xYBXlq1Ey1rYlR8LBqqB
i05rqzH2q1kXFTfegOsyOvjjgJBcmZ4mo50ms3EYltnBmFSuT5S/+YfPWFmXIo5cYDyf97x5isoy
ETjXy4wIpc1vo1eyPEFO9aHmXmqauAeyzsGYnZf9BnV0AN1BIUPheYQHCD+5zyxVwnfXvrdSMQDD
mCsi4rmETEyaMv7XHZ9p3vimTlO0u5rBJfG5zcsi0KPhIPEtABq2bt9V+iN5+YdocAQ48NmHkF55
BEmwsYWoSU++kmNt5gE5lK4euFr8TWbt04Kz5pkx2GMBtqH2vbl9vTnDMkTfXWyp8Yr7xQGkloRf
KXyIUmBtP/pm5819hIuU92wtNhg2Mdjsgc8nHT+BfTUq4zuxbi2o3M8HJ45Rz0R8+9f8UMvR0sho
Ez+D30lU2P04uQ/KaLQ1V8jAlTGYfc67YBIRtqwLMo09QYlB3SkmmGsSg0P08VXsp36uq/BN1gxs
qzLvoo2djX+nxP5w7Ynkg3UOt8S/ac89MKU9MpD6g9ziECeT5n7Fk6M1upJeWA2CH9W8Ea8M9G3E
+RPYOhEJ0DaPownxqzd1ylTuqdyIVwFdV4AnCQvaa+26/j5FHS3DqtY1lWnLmz44gYZ1LJvODLFl
Et0cmA2GzUwZajsLicmjf/aNEhufCUSn9ICkvW3t9uHCDu2TSlkioTckCt/A7WMhS0P2niIUko3W
xpH9LJb0q0sxvrXRbV+VMwEWAOmvjBpwqR4mfhtUPV03PiwrY+9M8BpGVfSWWtiCIbj14XJYbrOw
4OiKw6CAiS+lz4GuqIXiR4Ht8tUOkpcwthpow5KSU7H4o/B6xld15HIo+xUzWt1xi08oBJzpBrfu
MfIoLmEZuYqnGhz8cwdaVt54ws2gf+rYk0cCqItG9T0sOcwAopa+nuhT2eLAV1Y8kQcFHdP9srzU
pVAaKrbgCI2JZla6Ei8Z8ivhRGwu9Qpv0NVZDTZHFzvoW3aCNzpS71aVvHHu/BaPA3+Q9eaUVkYM
Iujn97tnOPUY/lcZSg1NpSjdPDZPL8hLP66b9sYN2wRTaZSJE8rJzmt9XsBYlXy/afg3z3uGoZ4+
Kl8xC3bS2+yBIzFjrFIZMJlusu/iF/i40IruXCePVppEaFmjvjyklVfX4gBYS2dsofOakPaz5C+G
opWA++FnX0t/KuVKsWJpgDEWqyi5pMn1eRrHWWxQLyHwhGWsoZ0lkHo/kBE5ChY3cnXlMll4VJ1l
RObgWjr4vsIyTzT+Fc6pnTXtbmj5aCfMceBvQAXjeWWVKgwSVeA9n+QMVoSvZjB/OJJK4HXt3IZI
QN6SBDvFqhJdiNocLeZRUvQl2nsSuzw4AGbBPC5V4c0nRFArsMniEWTAS7I7kDCL6pKV1yFqTFJY
Q4ZUHaQN5kb6bG/VQjZLGeoaFzYRn3r43ZGunRhylnVni0Lw2FMlgyQYf27Na7AAqeVUxYkjfk/L
nTZ3wZ18o5cpo+6i6cU9jK9C+sk1LNtw6gzqFVW7Ra4RAXDfwyBhrfWXWe0bzQDGIrsiOpI0sUcc
ErWCC1umXPCCZCHeJGI294JRiCJ2cXC2R2UL6MmESNFfDcPhlW3zBBYH+FLSzMBI80bdRFfGbO5t
rFhMAvkfm+lOLBcOIlP+wdbWj1qNc6zOhKjunMY+c1/Xo/nNMUEzUuZ6fLx68G5aLB1Tjct0b3ce
/M/6QEyHQNH2i8oHWAKwVujuAIzA3/PiJfvlFuCb024Ejb0zjC/+StL2c68t/SPCA38/aLXSfS7i
gf3HwNlOLvXAXxv/Yv1os4yXBelDAUYTZoyFW2nnerdVg9xZUgEQbi8skWpdsfnpzDCNvLO4MA6w
d6ya860V7xSRb/ozFSnKO7KCulGHa9r2i65s2IpgvjeqMcXHiHER4SM4iLheXNtTQvBNgiziTyPs
hvl1nYyUAf2veMZ/E9THMyhN4nZVCTf7kXTEcFkSOe5jPLZkklTEIjt0mbz9elAjGLx/u36C/LYb
pvsDuwmrVdjr1fK/Fdfbkqx3M4an4a2Qpn00QrydSbmIXaitYia/ovRn5EradkZnloqkwb7087nR
ztWxZ4yAx+B26wsOQ3MxmRdKdZnY4ElimLe21u7AwWM9FdYZ/PbvrUFXSmnsQqr5BnsL/sBs+Yz6
oEJx0Qqd/HanGaPBWH/pHVkNRJADaeMYs/MZP4NbPic33OoScGb/rcFbSNGucKoeWTiCLNgJd0rD
eH9yPM2MogN9sIP0hzhXFNBr2HoYXFSLZtuofdt/L/aww4mQX1ugkoMjjWy+Z6FgqwFBsj9hVOEe
dt6mMgC+p/Ed2j/syxRrgDRcOpqkUKpXdApMEqjVM5x5IDdUFB51v2rYz+zLrarJcZQHEqZSYpHs
MKH0bmEcObzgdIdN7RXyaQZeaaj9wybYwXshVOx83rCUiHyUF7K5qwgZy2iLrns478pABB1WgYWF
uyhCkQXU46j8Jza5HyJ2mAeKXeCVj5x4bXVTWlGU0IdizXROwh9uKE/8xadWJmiThk2/W95bxN/u
HH5KpctG6vv0zG3gK4x85tHflrdnwlUHvgkRu57HHultUsSYk0B/s5iZ/NGNcG1ps7SV609m2lsA
CuCYIwnRLONVs+G9U3YZZR/Ly4s4WDbRzM/6F2lV2gN7Sa8yuC/8eX1djOE3czPPve6zGtErPYBM
oyuzsjqcYJxrB+cJPoDR0BC53NZ1Q4V5FgF98VJQCRZ3p1aiJpfkMVE+k+Gh62tz28aGvDkOo3gz
j2UEvDiKnNtM5/A9XSKNf7rYohSaxswZ8BXAj+skWQSWb5OIN8/AyeBKHSUC1uSYcbtd94G33YAP
mF3p3cYNIYFtVMvYt92/TX4bD/OU8pXuit+mniSCN1iggaU76WT82oOeFryuEAEwhGW2r0nKUgGg
z3i4IhBC+1mMXsWGrhCbtB6GFagm7zpuX1ydlIf5gF4bRvpPWc45KLioeYotdcX4x+N9s4xgAM8d
meG2Kc0dY9yDR8t60sDCFcSAVpASKG8aLbpwEJ7N9WyzDGRk/Jl52yPspxynZHYQsUt31ccOQuRr
FiUnVFMrk1ruKJwxHY/qCzwL1LzPGeCAN9YUzdd8cMT33tbPLT9l5S7m75IZeeMqY64Om1vD1VXm
Wzy6L0t4IxIM4Xtwsb5gtvet2dDOBnjUHbwfhsFtECfZa//EtTETYrAIsiP60HY6Hb6idW+t6X81
k0Go3AB4/iCG31h6O29rUPtOsd7qCiBKXpKz56biPGE92QaldAxmTSeqscPBOXMf/pEvRKaFNMes
Q4iG6inzZiczOZ3Tw0d/H+N+w6yK/ftd3Rz66stlhs0amOLTfOwD+Bfp0C1dCXlbdSN+w2ITwAda
BUTHO+Wnhq06ZNeZ34VbyNGMX5BAJuSpyDo1xwXIrK1qaCOHUx2piQBIG7Kln/y75NbcMXHnVfm3
/Ypg9v0/Ygmta9s20DKkm6/7dGUy9lUsYzH0yJs/GmbMAASR75mg07qe0PL0M1VuP4Qms2r3buBB
uUEXPonajY1ratOzEWEugJGyzkGiZqJa9H5BsYjGWylGalRKcz08DoCxaqWLhVkjI/Xbyx/Uk1Vn
Vry4lOEWrf5B5rOMAi84/gH3verpRgALtcIzxSmsV2wrvVZjr5Wz3v8iFj4ypP4vXzT2BrxJ5Vhe
48JiGUmx0/iTyWD8LLO6/Rr0/J5Fs9vpVxWpmQD55Ml+b/zubwO57K5Z5BGgfjiP/Qa3YG57uWas
JpK+M+Ufy4695euJpM6nxCyKwn2eXSkSzgYm4/KbJY6lX+v5qO7Nz0gzMM/6zL1tCWfsqNmTr3BB
1TaLSxPN7/+rZEGqD8wsheD3TogSb4fCpQmp2Qh8PYiPdTCSMciTSlX3TQDBjxh1aPxUT47Om1Z3
soXB+mj1sgweE1qoRv5dPCqI9J8G/tMX334zhtSeEjnfQfS2m44ZNS9sjaIwylqRX1nRQqD5md3D
c8FrzLKm/cGK3WJSjzgSrHOdEPQdYzbYiP0p3KGlktmFdRCA0iu6dXW1l7ALu4OMYIpG4P4lDtmI
Sgfug8Ag0epU3qqY/esGwqj7Wl/NpY9OlFzcCP4yP83Kry8HQ2AB06q15Ki2TCDKCL7NZoFBK+Vg
vT/kbmrJHjsqc/vPUcugAPeP5jBtsRkaQjP1xi02yRuwyENmd5IIKU6zRJyUfIY+P7Q9EEUtqPkn
YRv9s+q0OfNeNMjNITjgncehJA/ow0x0rW7lHM0VOzAG5swVibF0Y1xDbMwvlyRQoiH2PaUeUjwA
BraUC0i0nOztwq8Y8RAt7eCI5ZOlxd87dXDe4m+fSYNz8JrLURmW2Auq8x32qJjgGGyMD4Kc666p
Sr9brGrQpQjk5nwrm6Ru9PGgA3/GfBkjTacuR7tslxS23YXZX9+EJfoO8UZFKUroIGiRjD5Q+kmS
Tj2pz00hmE3iDkZT612LXBPz1IB4ViaiTY3G4BC4yewtiuaWnJZck9dTEceSqdi19qHMpbpLGKH3
k3HW2Ckvyci6UCdAb2PNIGLuv0626yUVGVppGpQQWt0rHzF6h+grg74H3NO/hFSJ922tDAoYDprH
45EAqDd8GxOD5Zw8QV7BCy8VrrKnv7jDDiY36maHfBdn5ExFRC875HFBxc2FMH52+lyKRgngDvcz
v39ji8DGr7SZeP4xpS4ss/fmjMG/Up1BStgPrgccVyHYHsyxpAVmXRvO7i/l93OuMBM3WLTADBLa
hwWV5G/3xs2Tqz/Si3lsVSnCG+Bw2SilH13+3f33BHxiLwey/bNCvmehGTBlG7mC+CxYbE5CPPiU
Jc6tF2y02K5FlLZXAetug9jpxemBuJGRoetsWLNrje+GTi4Nf9patsgiwk5dzSFEeDP2GoaFA+jo
gx1WO4DmilOwv/aGxaQAkhBOVmxxKjDgXRUzlbJNJ7OX3ishV361lW3VK6n/WRAYE2u6EKmS+X1c
cXNVHdgKZMxgjSYPlq8sv6RUoeYCUPiFqYgUFE8wxiFuViAqyh886GC8XflL1AY3pH4OIGur6jvX
DMj33H4WybrGUqMf+tNQ7YfYf+niKd6J7ZypFqY2CX985sHDX6IBYiKnaQ+ZXJp9JuPf3kdld0Al
hxv4ufuDtcJo1A7GPhjFWVPy8FEwAZWqPybPRMAAwUss2nEcGg4Axew9aWc16D2kV50t7ILn6x2P
r8fm9L0+MCWSYgbq1EENdoZoE+LRoaySt9TqVn1YooDpFb54J5z3IqJSFRZ5OsoytqxSgzqNDJZl
R5oqtTuw0Wxk3KRgYAlqpcTwKFNlBrXa1eI+lY02VZzaf/4WcowHOBhM259B7NPQWX8yaQ0SVOIQ
oDNkTN9Rw3YbaaL9nziNt3DzJcBu2zW4+fHnFajgiGmTQe7ZeNCvLjVqxoTGgKVzlE7H9E+9lLUP
CX47BoqYYLt0B3aflnunxHxZ+U0c5oY6h+t865VQbHGmpmgW0xGaPGbsXaZQ6xYtO6sjmvHXSc1I
3tcmAd0SmoJyhG0Wvbqq88IQre3+L6shi8uT1Rh9F2c3X+1u2vg1uwgFDTghRkOePN6Jq3LWkg4M
PUQzLDUWNSclN+rUsznYaqCpHJxVoMlvAwINvurXDLtHE7WPVYVP33+ky+I7YRQ6/8nspaMDjX50
eM11UabqvegsuOgWhtUPsG0uvVRoGC9VWc2ffEU+BbnQd8EDO4w7Kmzti72DAFXxCKcZiRaAdmFb
gnMrio3T/I8INinNrYzTDsJy3vUFoB9E9vg6Cr5iKztR1GPtBWT/aKBlNix0P2AVVBFV+nWpgo2h
LDKruYETBv1kw+20/F7edRphuBFADyoK1lj2Y80LYTKrprqPEO7KeQk4z13VLjQf9RyWAif++T7a
9vb4KhznR3NtSCaIKGTm5nbyqkTvJin9sITQ7OOM0dJnIVlKtMMkW0Cbg/vNg9OAb/bF+HBl9bHw
WkhqYjYUyQBVSUGhh0JbqDfIBKowOqxNJqXLlfNgjP0gdZoToSDXjftLLTPG68VTYsNb0dptI5y+
cGbvBJxMctBxqqn9fCFwbr4XnwlqN+mUiKBENv9s/TZO/fETnJ8tn1r/ASIuYmn90+UO0gKUxbCe
dJsV79bFjCkJE7Nsl+D8J62jjPv4NbfC/U9FVc4WPpD0Uciu3+dO0Kp37fMJ4yPcv+90RScxXjOD
ueD4VqtOzrepchexMHXW0FFhIsBlH5CexoN3GCdXSyVI+ZW3xhhubsQGQhV74lo+t9jFk8UHCn3g
ybWBAg6hHbFhpeZNO10MaFGCegPJDgO/IH98TyTqtlIj4mNNzntz8TJ7Wcuuka1xwsi5B8q+ITOm
h6bAP/i8rFLrsAfH50JbDYzujfHmYUG4iGbz67cyzvKFtIzY4a/SYXwdjFGMyTZT0xoyLfhGoWqz
0QpiaE5g4SAVhhxAgEjBHBwA2zuR5vyfIQD6g9e//SiCNgIt71hQEFSEyntcq6XkB2sqEREx5Bb8
87OgncnJBkr1MbRBazms/bQ2JIOjFct/L1PI94UY+MmjgourabuJI7KFhwyDI1qXhGuDMVbFKC7b
6wtC4VOSEmImg3NLyagoJA9utmJm2jm7ZuMx9slmlHC6/eo92fGfEx7kXR3TjEOr9BRO7Kxa1SlM
c5Js4ju7/n3UvhOwhGSWq+8jKLcRVlgpkR/NXqd85kIHxxEV73N0zOR9HpuwiYt/RMTjer6u4t17
XZY5nt5rBHbYRwgRX9oGvenD3+bla3WriRpKR+dQLKK1yCNzqzNr8Ld1eqVJX5WQCGxW91fom8Zr
mImNGXdCSV9ZZxuxadlk91abY5PTY7oye50B4WHPGaEiUEqHqwoVJFucSEG17vKSnVbvXbGssEoo
6yEg21kgOjsaJ2Ggr4i+NEZJwstg3yv9IZ3CWp1bykoO14RoIZloX1p85L1TjrRwct+Rpm1cBu9C
sGtkfGG6aRqGMCw2pSOUvF5bvdJT6APjUjyi7ET3sc3/yyMYw+YccCIFHb03ESpAIwgz8NuRWzFX
zERPVHFI3D8Bta9584iUKEt+HllZ4HNUzFRrz+GTF6yjBe0Us+u5xRRrZQ4MA40Ma+5CCbpISkVV
6pvCiEnCDakcb8SCvecYqQ95X6BjIkUxbKXGqf6BIvRLGcKB86KNZM8TULt+6HFrUWBzRuRde6Cx
pmej9k7eXLVW3RM1uqcLlPr5W8zb84yqSlOa1A0AJ52YIczFIe1SRZE9WCOqfbfM1Zmgulk8djAf
gUIyKv6/k0G2SzsJUKb3cPpvVWy9E+is7dsFBbPeP4x6H1r22HhoXhk9ogYSYPCv4+mJ4j4vWU1Y
ig9/tpgFc6tsy5Y7mpTJMFz0FLTPxaylnKri6GEhkQ2aM7AxNbGDnHmT7iwB9kN5RxYULD8GH81B
qBVpeQjIuagm9+E17EqoXL0peCQwo/ge6fCJr3OqtAF1e4txTxZo7wwmI3AQE5yYJd2viPCi0yzO
OgU7SDCBuOQ5EKb6sHXitL1D6e3q1Fw0/AUEthD6XcGjuBylJpD1x56kQNhwBWw5aPKiFCJw5dTN
CyDx5of23HdogOw+0HDDA481Ao4NjXqKCgJM7KoQixxruL6Gar+tUz0L9APgWy+KTnMGxRgiIJGM
OfqEmMFiNtJsYKcLJueTrjq787/Ydd/PAWeDkGwNmCR/N1q+SzcOZQfNMbsVKJYpVN4Lqj/xqeaJ
KZ4W6LmzB15tJ02zWtYDII9YaRyjvjnBIYmivC8Hf8uIZWOQY4NlZ+d7NlDR0xl7jvImoHbLnXIc
U7fqVZRKfcuvAEz70WCeqHn4W1w7W3Pxo13NJ76yNN1eBXMk8TlLOUSiJlGeWaZNwc4/rkNI7D33
AgS6rRgWXGDMyUFcyJPjwt6kkcRoIKTFh6XDzoF+Tt2EEZ8FxIaI2VuNAbkctapYa8E9Q4kxIMZl
x3UlVJSUkcJAx38NXVVeWPaQ69Gqs7ovNfnem1dYJ/G2tzVoJVETIM00csftqNAkaOs/+rD0VopB
B8zGU5RSc5xtbcGV+AwmbVv0Hi+6a3taU9dsUEGadojmElaUt+9GivFDBAg4JkYrN33DVBd0EjJt
pN7xBija0qvb88dl/8V0NaR8k1WLgnhBUd9hlzNvqtbO/sfTEXYbLy221/2TPhbItAwiOrPnKU9v
f67O3RR5d8UBHNpy9mASllSA8Pk6BnoFwKC2OWouZoKDhyHymNxGDxdqWDtGbwkh5j1pRGU7I/bo
vWu3Rt3nFVF3HdskgkigJyIA5jMEzJNaDxft2WmZXKInnYPuSZV20wOaGucFuTQPV2qOwM23PWBe
NaWY/77kj2cYAFQsHLfVFcyP59TEHCuR48oQaRADvcFyEocJH2Zt0NU5wm4W9B45Qk+nv5KIQxdq
/aqU3kbWQsONPGoBATof7amO2tFrPExb2N9k+9T3tcDlym4t9ZWhZVxkAHYjl7O0co0c/EAEHWym
TPAXyy8/WVbTR2K7Zg2GQEQyjD3TM2CdmPo0OMuFpLtMfEB0vFKsRB1isr4oT/TwPU2Ibrf4+DB1
31way4hLg9lThXd0Xfs5tKX+xfFm1nEtWfXT4Jc97xp7prO8p0SaOp3yptnr8C041VKq0adnIXqi
YLMNiJJDyXIlORBrlQhaoN9GM1oaLm63pnkFEz0QKCDsjAEsKVGlm96NcIdoIEIL2RfwcgrScous
sO2pzNkZ8DYoa3pt4XJ73fOQ/p8WZMyFtz047Y08cUM+dIlUAfZULlmx+DXQ9WIdJNJJpizi/+iz
QBwP30jJLcn2ZK/R0wwMbqf0F5jeqFIFpk+qWn6Wm/DkKWBH4PgnrREmn/ItoxexeYao3Em3XzI/
XbKHhm8esJcBFlN43dC33rGnL6Lpw+u0Dkbpq1rYvnynJpsASpSbXIaGNnMG3ViuFjk8cHkIg0nU
RWO5ZSKid9ChpImjqc0jQqDdrDyiJc4sT5UYsCiaLviZdUKU/Jxo2kUMb3V1/LRvKKDKmvWCvlE1
VFl77z82PDHG6G1lFNAP1d8TizU5XPNiFAy4htTl4OoWqLdCbANuhm9hNFhQ0M8vmpGOsNBdTqlC
0LKpbajpdZfFd/Ef3Hl+dj+YK35qYS4fnq4JbHZ/k/m6/poHSOFKiDYLOQaoF5oOCNUURSLwcw73
gK+F4wqGEKhQtKDdIxIeUsoADaV4P+YPHLJJtRQn9yLWPOpNaRFrjaxXCB74CKUXrDCKRHaCS9VE
K5A0gDCP8Vixulv+s+AaZIap77PWJTZtLYM0BR4A0HkcvZ4eTX840+UU1Fz9GdHcvBqn6iW/ZYxd
HeOWKR/4iX1QDi8AMmc2kvFOPjw72rGU8HRwhF2dESUhv6Mxehsmi5gwTljpgNG9EWMXujQag4jM
fRnhlNh/gqeWYz56A2nPtBj0XIRB2QGYAFE3Ue5Fld+66erz6wx7sDHZ2tqOyKi0EUMhiZtqEONY
Mwl8EzB+9+F5sXOEQuTWUNJchpGiKC2BkaUZIW+sejGBeYMCxP2WVTKtC+mTzd0zLdkSZ3SiIDPl
k0geIysxrDvowGzP+ufLBHjfp5ZM36lWbAeE8gbIw7NcBCk8eV1xe3Mqirz/Z22v03h55EvwuDew
7dOFykkt0VhPAtKZDtCgYbKeFhTv5J39V7Z9zL8hwXv86f6ksQbFqnGDuaktIH4k83KARvt3d3Cm
tn8e1MN1Q6d9kZVPUlwKZE1o9QEzyldaKSpUV336Gu1GRalPXbKkmK9Eg0n7pqTMaKmk5vf5YivK
gd7IWCzQvlUoNqUUPT65QLtXTxRtA/E/PNZkg/bV6lE041slem4AYBW+jlzLQmSQqWBlZfkGFvRX
piUT4cihqvUTa0qHQpvcxquDOBerFqSYNe2xNcbwY36Okyp5omMEwzcTzIzKqdZiK7kcgQKDNXxb
wLORw9EQkoMsRh0s//6lb2i+AppXduVlLOQEuXxMXhT+NxRBGYhFXdPuH5umIBmBvF5FesLSxhU7
rVLZCTh14dipdq75ULyzDIdzDGPlarH0zW+p83LtpVQwa6fX0oZDlYO/YNSZV1NRsz+L1wTM/a04
FYxQb5eTYH861NGBV+fuS7d2eb5vpio/pQXTaHh00ES5XHJccQT0t8ZUCH1yPHnJy5fahhXYWG9C
hh+C5efsAvIMxFqpuIETiXLOIkfuJzXln2Ng47Ry9cPstVZc5sL2r7j4m/TwkIA55sNV6/fimcUL
HLzO+PkNAPRRz2nqBTMPuAoXPtv6kAfDI54ZtWvvghqMgObicswULwAyfA2tnrb8A0YnCcDRyrpF
1sJgqPGyzmdnFFFA4VTxcdRD+pQ8jIj524R7rjF/beG3WGy8U3x0sHQCSH1y00uCKJOGATvz/Vvw
x5uxeeq7Mv7Peo8Zs01cMKMV2p+e9mzAb4sOHJK38VLEs3E6cI/8nKOlPfyt+PbjFC05TpvT/5O1
ZymNisH1226DfjyfIwMfwmIvPz52tjmu86+Hw7HYPqEVFJeSmbgD8yernl0jMnIgTLRg4BBFv96l
bIE+VvCW7JtH14qpS+5ROvxbNfIWhNc5ldTsLwDNQ2IQmHSDjhkKIa8Ekeok5p/gPLOya/4K8MP2
uMh7htYkJXfg1lvsQ1twwJPty+s2h3ahrxEQbYl2T0SnQuo6zOQVtjo/slOY8fBRzd1+u2DySJSI
GW4q/earlHzC717irMWL4A2O3NcvFg6cqONeEoxmGIHMbxBS5JzZ8QXMe3JN5bKaHzD60mnsthRU
Dh3r+SkRJ1SfantM5xrD3SovaNb1Gfmb9pkIQHf8UT7yaPVN/mPJ565ZripoO8lPiGftKfur6GDC
c4K8a0sPijnDDi3pyk80yxZmVO6GPrRPUgUmeeqiIHMoqahn3DqCx/dZwzidQq7t4wrB7uOV4SYN
U27B6+m5NTGmB6+WYck/sZTISLpkFD3vLKiO+fcVDFbsrFG4gZgQZ6e48Uix98MVCZzJnVa5w5PA
mhiZUhQVWaY7punE8x9qDEEFwVLc9BDM766lpewU80zPwdUJ8MjTIbY5XFtJEjpLJp8LCBddpEx6
dOxR8o/tecVvO6yGVm7TptuREuXXqgNFQQ2rtLCU934ihxoeF7TReWvlE1igaOLwPxOE1x1L6Ugs
ym8JXq6GFWf7PfOD0Dov2iCB8X0d81wFkxwY6qHdXriOQrzTyISUOiyf0tD5K9joY5RQG0+5qqbY
W25yjS7fdQic8GeNez4RNocJcr74jggh2lx0W+OAmVL083nLc5AXEtmK9zR2DCxdMjLLYthAQPX4
P0DxSoL1YPW8YgOEBC2styRwx04FWc/nOCSBi7Giwn3X4cOQD3VqyYXblLnDkp8Js4MEd07zfmaY
ljN9oeHcMnHXFtkNkNRS7kHgf5CazPKwS8DeMFbjBfegDRGSmFWZmdAMasaJRZSPElE3etjxgfDa
B/Fvh/KiBsEK1Jq7wYSRre7I+c6MZsVuKfEmcNhH/Z1J0nK9BWFUIGY+7kPnEAqbqxhQ9iOYZuq/
6u7E8DOpk7p7ft/DPglO83NmeDVih8aJN1kyKMhUAKRmtlHcrnfSMugyV8Y1IwLYPHYdEAd0GRxF
QXgGAzWwjbL5Tu4cxtvqwkGjIhtAV5pecURDeQOVNoBmaoJPbYXQjO0APSo0+2J9g7U21GOi74O3
aGdeJC7pB45XtYRAK8ekfcSfWeP8GoVJHl78nL2NjgASlzfIKTYKqYaczxn6g/skdKfxNWs8HaSV
oa8kiqmSRk08iZl6UfJ2vrseS+4DY2nm2q4Czdx2XSSRP8AFVp2H3WqIwwTvmtZFhY653RwQtUFR
a0A4vJYSVWn1W0q7jrK8bmoeoqbTzwr58B83lPUPTFlLfQtxfw6PNATMehC9bX4aniraQUjVqPCk
s2hzLwwgck6Iuisblin3tvMGJMm3F83pe0hlxPUQd77wg+Cn09cbf6u8Vl6x8OO8y0cJfpsvV7Wz
VfsRn17+lDJSZuoK1u+WQv6TiAXyH5+p+F1U07hXFN9OOAnSy2g+YiNC2XorgAM5iSU3HT6v3tio
25ebes6Yh45kGK0a8MdhCGAPrmrkEt/FlyUIXSSO8GY5cr0MZWun5pTwZkdzcpF8ZMHt7SDZTYyu
AjGkr4ALLvwFClGILRuNwXDEYWQRbvdsFQQO3HaWkC/LJxhG7rmOIUwNlfdE3X8PqXQxj9XhqCa6
Rgv1D1NcHJuUyBXarnjOfWP8lOtL9j6P668oAmHXdW3MD7l0x/rCinkEG3T6c9Ve0m7DjH8dbRcF
Niui3pvFNayWXNxZjHjo/jkzVfDHXwQDWqRiS99oByjwX6DyDtoHR9jw/CwwNUzep/4Jw2pjrpTJ
g4vCg/6esuSS1+4h/7PhwelnddYqwxJNH3q2o28TKI8NR5gBcTl6ScI65ppkdrBUZooXG/m36zA1
EI9CIe7EI9fKpSNgUhbn0cw12BNB1BBgHArALjmLbGYPiI06xxeyeRQEe4qF3ca5X16ExXNiWOH1
0b3oGfiNL27tyie+rHJ3nbferEoM49kfn4GWPhe51Gqd5rw8SsvMUE3R0lQ+P8kzCWqaO8kleISJ
vOVhnTZtoWZOh7sFAWgZIvTIAQ/mqsJk6EMX66HzFYkCf75ib97rfQjkw5NthTO8vakuFrxkWA/p
sswHw3BBHG1CnkR4XcaI3Q205H5y0eVzAhQln5ShyUMj5ajniooj7ySXHwMYdmugxmhHkdnskHzC
P0MpdKwyKOX1EGbSAuJvmbegRk+UaHG8cbMPorFkQZvLZRX38MwLzTGIHX1fpyI3mwbZhDZpCkHf
DMEMuctkYZKFJNzbc4PmKjWrqxqP1Q6rhfbnSz8d77WF/7+7utF0D0am4yMnxUGc8GURmgGScrH8
o9Ocw+IgOyIg0xbqzYHPhkBSwdga/eiSjBW3wsysYSdhf0P9s8UsDRlrOl8FALvqgc/MkJfpIZPc
yxvfzy3zZ9+lqKUG9uHM/E2D+F6N+pZ6KCfYvcy3KXqkW0QEQNftdGzx76gmMZBa3idxoSHb/kDV
NiEo+KPiw6k4e8OKGeg6S+BQOwsuafB0P7gXWhIpXXmyvNAIxpYpWgJwk7+iP1FD6YFxJhLoXNwd
dYvWmd1yykkHveb+3RCXh498CXLV8Clhh2ggXJuVulQzT7WSLsNU7ho9vuQ0y3KlUrZO2tI4pRbr
IpuDtJurS1ArJ0utnwdzqnIXgO0zULwdEI8sdADwi2AgKvbf2QUv8ARYnokCcKMOfo1jLhxns8nP
e+fE8T/0jX857waG/0sC8qPNzxkxhPzv4x5lFao+oGDtdp/EHprKRtwv2KMBOzJ5ws9qpR9Y9pCu
Ak0vGGTjX4/On5zwqYz/Vkg8Q6zG/fTPeCvPQz0xOFCavspP0eaYDLjHeevIS+EfVfd7vkmYd2/C
NpZ+fqgQC9XXJdg4C3jKNLOGQ8Xbhs8P2dHfZD+ge6JjiVN9eEhj0QOGE0V80zMkZr1lTsvGe5Qs
qdf730w/4iqaf+Ww02pbTi028imUCeJWdeHImcxeElsh47Paq6jTsbm8ho0xGAtCPr3gTFUlfVO2
xSKtKXpzrURo8WNfg1xkgm4ECPI4DRIoXwufCk1ju44DNNTGTK+rGx8wnIAdmriAAaUMrSvgF6dw
K+Q58fHvw0L/fkT8tsHzFsluxJm/avSdy9FY155qAlSqm5TIBN0OHgMg0nn031PBpHwUayUUo6Pb
X8dLybgLeclRuZvwdwyyY2U2YRH+9nQIwVyn5GckCiRWFng8UG8I/YRW6uXBpoAVKzdOGMkQTobK
eVjJNBJXRZVXEwJ4TA+ZqYFv/XpDNfQKTvqECwfgqxrB0QHl+/egMLuSKyh7OImGsqZHOIfavIZ0
6EzKJPBcELtJmzi2mSiDwYzwThM4mCIOEI0Sl809DvFKKzQz3FSudlrqAA/L+6CjiNPUm3HyDA0N
0urlywRaFVJDXciIMsRMJoh1d+pbY4cu+QJ6u0tQkEKKrqo2ueDilUxCoBxqfQZtN1bUWxkzmRFU
4TYI3n5HsPG+I+GyOlFwqqWq6zlQ3TzWl3lgta34mjt4VmyjbaP6J6ArBvzwIvuwJNyxb515i2Rg
adCkLO1qipxLbp6uVpZ3WNjDqhyqCeO3Z88ikIWfaSLTc6qswZWsnllZIoECg829V6BfVxiGDDST
mYWHGL9s17Esv0m7e/g1RiERN0d0rh/Hftp3MHwkFrTaFCTC/bSYJNcVgWM8rrHUzTmUAnsVAtuA
Lz1p9G9iihsuvJAZP/r0gHpVp6xoO2SeR4XY4xUeyXMxbNmDmyyQJH8+ClOCp8gChWlgzZo+o0Dy
Kk8n/9vsZLThMwiVX7hPWCjtmL0KntPma1LmOpZz9EzebVfZoxLYVcwrh4/xKvYjHzYpyRB9ospV
mLmiiW2/OQibnDd6Spy5AYY8FPtOw/4klu1porQ0L6JsWbFSUT+OcMhckDfjp/zF6gF208mkkX82
VqkNJNRFmMXRQALQeGMe5wPDgLI2JlHk67kCVyXHGn/Sy9/YZmNnCAhM04voRHQzGjEalAur3Kcy
sLqqtw5fKGRrdwszHQTMtL7qORQL9Tu7J0lci1Vc+hYNzL98O8Fjc5ScNdKBpjIdHMs/mAfdGbRv
I/RYaU1xlVk+duRCfJAKcatqCodImczTYFolmBIjynqwmsxVNdQsRFZCRoAgC5m/ZMmIT6nnl36c
3GoMcrf3KfcCVmH0pOxy/7vHdPLAhLL436iY6VAePcRfU/IocE/j5sjt9sep8YzzyIo4B8rWoTzD
Eg5oAWBECM9fr3DpxNuQXwqdYrJaX8UbL1lWyCH5SxnSSUKisDo3uqIW7T+kgj0eIKuTbGQnfIZA
W+JOJcf64duEsOhsuYWfMv6Fqx+kvt2nkFnS1P15kPXJmHnl4Es9/x6oeo/oN7WxDA/YU2oAmJGi
N25Cob6X/zqWtXOnhFIjgyX/0yZmIsIJ3gn3awrJ6D21Gmqvi1l54X5zKU7bCBza3LlXh4Lt3kUO
28oUSKU6eLEfm/IX+sruHS1ufhst/lAOalyW/sNKwfwT1Nr+tYYKHyCvRa4mgX7+68tI9Ud0uGHg
3cYcP8F27+oG78V41VnI42IdHBD+/3iHivUflUVOBez69hIgww76gsh0df1/9BlJIPSILpp7NgAp
JuJhO57Y4hArfM9EMrPLCdp2zAod88gFSYP/9wfMVt0UbodHFKkJ8pjnOvr4kKfEXML68ui3Skyp
dXnE2tmekPHD+4bAP/xOGsUEEHsB58N1K6O6T9+2R1bFoljINuiDwQvxrnyy86fIkhbpMSmwdA/x
+fCdlwYgxH1vag0RRNhjF55x5gsWgPrIdqtEeVsEpUJNKMketNq68wU76XGUBZjql2dW2/HeTZc6
QMpM0cMKtMDBTgW4ltIrMbQCaRS01pXpwRSYFZua1b8+DsVobGbjdR1rznrgGFLAKffAmMu7ICw+
R8gZuaSsz5e2I3dyeaiNCGQscscBogveeFmx2g8PnFx1F6wpGxkQcS8Ml6fbCbKlWPTUD0K5HuPe
MZxBt4OIx/3qKRrRDWjhbjLER4ALOGxsxyhv7g9qOmM3l1V82sFWTgPjmxT01+Xc30fboH/xTSIA
7fiBTbWpE870480xPasnLodjqb299s+kLcWiG/yAYRT37m3aYRJUdrRm/PpwkQRZOHorIOyFUfCd
1ffxDYXozfWSUUhgittTTmcTzgK705n2njwF1tmQguxLhB5hX8SZzbePVqiMACzI0iFwLHezz+CT
btwpACaVkauKuZ1gOGVqZamLy16mBfkmQsmyAOb7gy/DIdTeNDLxNDpOwoOoLOb5xjH3c8NzU4o3
0fnuPosjCFitedGI9dvQifdjziGNQ5jCmbqdM7N+TP31A6ikCJ992bgUuoWv13KmzcLLyaZYBbVl
UDlvL2PO9NUZS1gxVK4tIPQ0S89Za82epypVHCSpwDXq8e2xFMeKVTOF0YxANbFozY+ullNl1qgB
1BOfgaVw82bH/l/49VaSSQ37QQwyG5jfDROh6ZtlxeYjjHGIX9DNjsHAY14/FJcv+uCcMAogjk3s
RbIKFwfwBvNg1Hw1DmIO14vZWSFz0aJhUHWMU8iStYk8i2w6RdF882v1uSwMPJBGwDuKKT6lDbRc
1NbROdjwf/n1Z0bAtxeoV75ndwoBBgxn0ZxJIJ4QXDFAiBbqLU06x/xrVezAdZX4v7dQby8AufSN
JzuYY+HVT+arze5EczZUnJ5aru5Fq3BED61SVtSp2w6C/1wJJoWaIK9FsVCPf4t/QUjxLa1rtkWc
tMugR5ahtMmr7gOVZrqpTZaA6fpNC8dHwE4fle+eTUi3peMPw6TlR6FJGYTlE8WQ9OAGGBknUxNR
HFr+FUgC/4OCJxIiSfm2VhdUMyMc1o46xn8iMi4nqK9pYYyh4Jy34iS9Wcm17zuRDQRLhnqeFUCx
fM6pGX0Tz2UCdMb4aYdLoVOULUNujtkVeI9BYzcagS7YvSvRp9Cjx4bQImpwn61vMyaoAMhZA11g
zgyqHL7gZnMDcygSsGJoDJow2R7DE1FfSvIw6BId08pYZAiQJqk3uo0dk3onS9sCjHFNV00Qougz
uc3/MGCJqwIO7Du1/2cQvnvNFb9LeBBpyfjNW2trzXhG8jVTY3tnEKqC/0BNI6vOBJmh2yxo37Yz
xQqABbUzPJkElKqLertoEMVmp8v0HPsAnGp/dFF5LSdhKLn987DMK/iVTPpohYt8qpFNux+KyTug
nyFnYtHmJ+nVPKd0/YA9JDplKswBxkMQP5GKfJpseRMltACTYNXBPRlaLrTeVtxwjBAp/AXcf6tl
aNfhUG/3SW1RlLeTA1M15rK/FdMXv47hwuJn7qxxdqadbFr+3mKpMnWLtQ981k3hIs1vi5CefhzX
TWW0Z106uLHM2fp0hiQGuEejFiK0UgAZrZtnSgqRmZM5c3sjqROsg3OT/9qosVsgbbv3Q5jSoC1h
nkUhwhh3REI051Kbf5Fs2x6Em4N7StKs6sPiWaEc6OC3PGmXsLhz02xRaPFciXDz/N96STdJvlJA
yVyyq2krfmGM35lDn1GSC7tWY9KdLMfKzvJvJONhmtPU2867CcE5Ok5rnj65HBXAFEuludXieXRJ
OeE4Imk1QTXV2TY3P5gpQgoQQDpEDtZhacxsb7Gm0NBvaZui0wh6OU5ngJXPA60Cc+Us4lMuZEHY
XB/IXh+gq0+kc3PFOFUCAHS+f1p4knsL+tL1w3cdh48OPn8AyD3kQfPoiOmx275LpxpCOujy5QcJ
iLZ80GyQsuvrtvUv1S0aJAzad+tjclpQfm8QYWcEjEKpABcHDovbbtgYyJusrsE3Jh17QGTtbKks
a+VHPbYHatadfw4uG7TDxl+ezag3UO4qvAd2I4AEW1NuesngFmlzr2Pejq5iK+YZiLimfqu0aTI7
xvRgu+ZdpwS+zH2URvW3Y2gnq950YuoblE6uzQ5Mv4n2DSYxn8SwRCaoklDU68OigkyybBTGEd8g
+CxwFgJjqQDf8dnAwz7wL15WqwmY/0R5lD7bm3miszkI0Whw1qsfLDZKH0j3qXci6tMfxHKG0qnn
F1vWsEyJmzbvnS08KLl+W7lfzoa3TtxD6jvQl8gJQ3KtyHQLUMQ347D587nZZfOza2pZ32wlBfby
Vrm9MxBCbnXbnpM/dz2waXkLjpde7uaAApw9cDUUSrxsTEK3RP5TVn2jkfysg9RXtwL4tjAX0rP9
pKL3sWF4c+jio6A81sOJ1JZLvmWtbkfAvXjF4rHLctEeGP3lm0RqnTS3C1DGh4TRDNfYXJYk0/Au
zg0mLtLXzVfjhO4i1Kj7XtYfqrhd6yWnUEOLkpyDITCHqo0yomMkXb10bucukaJz8uVIT+5hI8EI
SeIAV8zcAALkcLKe1pTsUcUh7L4aIp8Bh4PZLj1d+1rGfkHuuPKY4oHiOfgyyu9tqhPquJkX2MxR
XfiE7AIggvT3YG2B7pjAKUfi/tTll7mXalMNW9B7/A8Wa24+R2znAVLi07NtaVr1jOHXgZBfB8Mo
tPCrRWNzUjMwpQaIs5eQcMa/dHQ+9b2AU3YTYJmY83Ax6C1N/zPdgpOW+1TVnCdQtvsOrzZMQopa
2aiiHrk+rCsfEBZXo2Kv4aBlVySEbozLZqfPp+MW6HBMHy2GxGGO97uBqXbeIyhvuC9WrXc+fqDx
wAXORVhJLyE69rVhtVCfbC6G5SqWUn6sZACXFR3ZZUdEdTi601k6RDY3ohECwhwrSYKOs0UJ4vb6
PmL6i1DB8tx2Nn/oPp2yHp/EhBy1NZn2G7o3UlMh6nSQFsgkcptoK3a+IBzjbRT8kbo7WM9ViTOc
757NB+o76FJ+5aEInhWuqswsmsW9pg5zIt7A2yeMUQmMH6mfik/vw/gic3eTY3QTwV9E2nGG4LDL
wSB1qoEEyhChegncNeNRy9iC+KinRMSn6NVsW91MqF5uX6qjxYL/kdMuEJkpT/L4b5O2V+fyCs+J
SIdZ3h1dkrEp3CfU5p8K8iubcVqMQNHotRbA5TYm+ALPGei0R3/Gh0RYDVvl9g9kCXfS0MwAjg6P
/EV3kk9oI/nu67oiTe15ugoo4xezsoCLHtq6ySVOvbcQrL1g2YMdmFhEjhfxQUi4i/+qe5BZftWg
XO09vhFFFBf/OAg0L2WYxBfU0kRJlS5k7pBT2pgVKBRjG/ZbNGblsVqozjYXR1v3w/jkOM5h3S16
cw4KY/wv8PMQXV2o1gAStsuGR6l/u06Y1sT4xov6BbtCvRjAjA1haceJFsQqIOUVHJK81u/5dioB
qliZn+MYF5Zk5qnoicc2+NVeWGiYLgepYRATpRh9D9usB3qM0FdeMYNtcW05ZjK2j0V2wPugrJVO
eNRMBxxH0f6POwA6OuTx/hxUHdVkwkxnHsXpJ8SKdcxRHoAc3WHsvSYFBCwasf4EXrs+CXE1nuhv
g06X8BZXJ+Wm+hwK81SbXl2DWtFFhrnmYBAaSPeDkb19AsSsevwgimYADPRl34M73t9FLQ/2+ldn
H2i919xfFoBD02APDHqWP+mP/MWJDsx0VlvIaL/UmHwCM0OvaSZk4Nh+FDr5zlF/KfCvcNsu0zGT
p+4ytSfjy0L61Wo3VmKWUBPb6RUZYPuOn1kp2kL8zg5/34FeLbyxQJY1l+U0shp32TgcDIFh2xP2
teGzUUSMh+Xh7AlFkflOXCdaa+HWGr5ZGzd2zFj26QiECYuU41jOp/W2xYdIXnyCjZAEAtVbCuCo
h6LYo6j3AOv7ycZoeTl2ssfdk68/tDRIhXjpQ1+NCmM3LbMFxITw/FsPOKWlUnYDVCQ2WBBOAxdW
upagfzG83a+CcM+i2yI9SNqV0JCGVd+eLnt/wI3IuzVmSv36kZbsxmG5jNyKau+p0G+xT4fVExed
GS1XxIHpPLUrPHkaee3C5tI9xCpZEmXhRoFk33eGbfDe9ZOb8kNt2meKEcuTHspI0rfwUhmSCsnF
97WPLOUCrCfOTlMMNeAUyQGfVHCBOqc0PkITJAG+TJ9sViTcbqyiquRrOb2MrpLmP3omXhCRhjeh
kgYgbUvndgHqR1Jbj1xLhNYMO6xz/DLi562041M1lb4WhUo0DyX5KbHkQ5Nx4XF37P19SRFvc/gD
atQiuexC17CjkNl+q59yytyCNkj/B6Bz6WUCrBpVUSv+2fBohapPweocLgFB4Q9KU7qr6yC3oJdl
0zXNSxM6lDsnRx4HAWtDODl1ir5+k5yClPb6rryHD3xdrnMuaZ3/cPSSxIbDU1Q7unfou/En5apL
AJxJxq6gv6bT1btKG70nlXzSmR75OXe0EwE22OcBhcJodRZgrkqwundIH3qKXRpZFNHKBJYHXOGd
3rBtQX7/3IM3AIJ+mqIVZPIldCB9dvFFxly71DMlFKyHvCGKD2rdmOEy+gR8is1zE7RS7+EL4Xeb
yo9WaKG3e67oz+xhqMoZT+FYdU+28WDYFnykR6mjTPlYccsX8N3ZLQE0TFPgjtbbUhWbTbw3psLc
pt+Nd+EGmcWXSpQd065ZeBf+1VoBpHMPEZFrkq+gdmfD/HaeWrV6vaBySwxASEeyV9eSda0q8AWH
zlOZEQCynozyAuHslAtpn6BDmlW2zpsmjwmpMiqBLK8aftIKNTle9McOeo8LUTsoS4YT8Q0R5eej
L99uLEGI6Nw+lJQRxSenZRIj9L7dBm+AzC3ifJOpFHXQPZh3wvmdtWKKmAED+7QjY4U9s9kEH/A2
LJY4C365bohB2GGcPokTADf3mTVutypS5uPpKYe62BOswTJdrL+fCQx0NCqNDGTsEIc3vlvkf4hm
eNoUy6K/Hu0e31SHNO8x9ns0bj08yYiah8y4DnW2+EAb7f5moxh9lPn4W+WeiuyLftBLXYcDupht
eeVG1lJFtIO9K8ZoDRn8Cm2EUBbJ/rfj0R872PhTFfQR+zrn3VUOGZ1YuXSI3/qjd+H0wZupaWA4
3wRoVfcymGL6cZwr8K/jFbFTfVwcFmCHcT6SKj/C/5e3gwcPt0AlEwNAKye+B2HryDBIQuR2CPot
q+x75Btt6LCqbzJYu+Wz0+f5fs/H4obzbJ4DpD0VZRQKtXxfI5nBav2afW425MgRRQNzcNT09irm
6OKYKgv3w2w5ep8tjZjXSIFiOB0U+zrYnorDvxJhJmouM3U4L1FaxarS9y0o/losxwkBBeaOg0xK
rbIMbB7fsob9S8EMJ44Bi9TBNz1WBXmOdSw2Nthy6t5pLd9Jt9AOWpkAZxeAQ+DJkDtrR53HjXuf
DfTFqTaGWW6muEwdAyVPmgapdvF9jyhwu42OP/TrJZ63DUXxUVs//8vFlTEPxB3okOxXNpT0edsL
2Kqy2z21bD61PfLF8PEfE4CJZ9FuUJObgLbA2/5/uJ/or0HKNHUsQsg8WdsBZ4j4Ie6vo31MJOVG
+LwX7bO71jyYw6LQurfGCoBo6PQtTXZNTyrBCzxHLeSFGSk4YY1mhcAEYbXLPx5PIMXOyQ7znp2L
tlGs70GQH5Owfv8Y9OIUiCkYdO4McuQ39q6zR1vBi7EdZTQEins6IpqsF9t8CF3hmZDuyM6Or6Lo
B946ST2MeCEMVTegeSwV1+rTKSMH1aQKDj5Qh7fSPcHB+CIPNASRBSX05zfcdqwi8NXBBHAill73
RC+c3KHePNe4qAe5X6c+vsIhok5pW3GGz3r+j7VGt6rw+DejXlueLwBAeY+cHJXrHEFLmMVlZEQ0
9hPpwLKG9rbr2c9LaDTnRzIOrAhLwz9kIowHn+ZEcfPc+1mq/YeXzDTF/9er1QTmrITDG4R2ah2Q
ParApQHPrFYzWL72xCfoQWWsv+KhQX2HVD6PhJM892pNYvoifWCXOdcnHR0KxaEbT1rOCevwHplH
tfujjW87VIxOZTTmlGX4GWkXzPm1ek9RbIi0rDimMpm4yzdagQfjwwD66sGc8G8MZYxtc/bkupov
zroSN/lHIbck3oLmVbb4ZD8qG50dHyc9QhnAXvnsaaLsWVuoMC/CHd05z/5JiXpvVkz/MVZjQPjs
0zy8zJQ5cBYmVnZMs3JPxWb7WWuAUJoeV+VpBqVHwY0qf/JeTwAOdKKO5AGg8K0gLCEHUfzl+Pp7
v0gh7IacL+LCTKJm8NFM3CMwoY8g1cwItOUL+5uUdIPu4VvZoAyHcs57O/i1NJ7XDe26VncVOyph
RKFtK2v3PsXMNhXymB3yYd7uVurlE8AlL+t/7E/c8lLxSyHQfxjpCI5aHAc7gctp/cTI492gEtez
iFbIzKVots2gyz+lMi+xQWdbkTt6iRPGZVnDTh4QIIvZRLP34tRRfgIXCWl+YZT+SE+XWdYG8LwV
ERpN0TEBnHxdKiBP2BTiUYKer88wG//zFwqEWQb//bSeFspB33weWoI9xThSxCZVK2wu/6Rt4sgD
pu3B2NyQoEZzqJYHvHqn4FigKNiTqeZtuGKZ43QEtXDWtDM3+mGkAuHavHZPmUmwa+hb3CHJXz0e
N1RmJPw37o/t4hEsykFVx4v1BiU4xSYnfmQib/tL2QTj3aZcvdYG7eBpADlsoaNUXp5E2RxrHYUU
ebLhRuCVKNWi1bBWGJBi9Bo8qZug5SZv4BsYQQMPoK6DV/tgYVYN3OnqsM5ZsQjsbiP9GLZkmt9h
tGxztmoO5yA4BCp/y6Y05VGUpEiWDbQxPvDR4S9Uq/LM0s0A8oKb44khw9bL/vDJ0wwgPURgO0pm
V/DfLql35MFWUhL0SJ/L8OFb+iVXj7jhcSQrO4Tmv/AYqBniFmYO26+gDWUM4aG+VMbWVWwUXX9L
0m7ZAmdcFpkUiZJZezRQ9vf/5S/XEDiJRkMHWjzcVx5GCS/2Nk7+B7xu55MwMnBhY+qVNcJf5F3s
yO3zS07q6eC9pi0hRmR64mRsZEX6Mv4C5rzUseYfIHyuK3ZB0nqICcoOVtSPJm51tV9b7Sb0MVka
CMA3XCuF8uaxyQvg6Er/ooc+ntS4tw2Jh7RiPzpRSvmnLOEHI0Nn3Y0eQPtkIsqwBQGB1PHMBXAB
pP71EKDUD0QwjFYYDrEfWV9Qh51ZUGFc9CJDfjVhePWCQaDZVSlR+7aAoMEli0JJz72NBN/n33Do
kD3hiQFAivZu4RxD/BG2UO9Gwdl0zKQ+aW7dw2qn5veXHYfJMEoKxi5mbNNqMxPyIwg8Z3Lwauyn
/K8maaMdRDujuw5YUPg8tSKyDeWTdEMMCzcYkv6GXLyDPEMXM/JqFaKGlahrnnIBgFkkeL3dHAOK
+AU7YiH79tQLCBEJE0/L3so9bLVM/Bq2fiXqtl5JpbPc03cAep0AveDu87xsEZCoXp4azkrqMzXQ
X1eEPy/po7i4u9lRmL74g6dbLSVeH5xPo0z/QatB80ld+mPGlz/0KnEJGdap1xLxhQtn84TiZ3Nw
a7kGotaPXTUCo6E5laP4zPYJFCe4gclcAL6ErYCfRY6C+vk8AbDMUn8pUhvlKnFyv5ZDiGP6Txtq
Ta/E5UNq1+ctroFRZc8NDoGXIJJPxcW1FLQRQ3D/K7NNO5pY2eeC2ObCKGb6PVNp95xW1t3hPWht
CwwwH8seR7k66ICg8yEKadaKWDMx6tHZn14yAqt5fx7GxtoS2mnEaRtzWK9dARi5IWF8p70JSqKB
2SWuJZvWzjxJh1ThF+8crer5TCS8Q/vX5c0upMot8Jlnqnyj1FqYedIPyPJ9nlWpIU/dQU2Lh134
q/C+EIReec/QqkVxsRZurdQ+L6y+n7x4eo7Ik9nYmEbv4fc5ThJ9BSWI9cDMr3HrFLGUqUzr2adv
tX9rBUfBI9gnqyS2k2t777kNxMKmSH8DYm/HeWkBOURBmODwvYNI4nJkggaYIw/YL8KRX9B2I/wP
aumC1xH3KXPx5lJvg0lTCYS7UP0yYPJ0DpxPLjPDrKkAbjhTBV85i/sAFmagOVPaAqiRmfx+917x
3zf7YUPJLrkxD67R7uOnDb6mFsBZWTizuzrr/mer7kgBCqKFiEDtgPUw/Wt/qyG/JRXQTboL20bT
EjW4koPQaJmk14dyRar9+72CcVh7M5OGL80NKJgwQrXx4/QAaUX1hwJPJKG9Pjffk7BeaMKvKufk
n/iZoDcAEdaXnsBtVDP2FHTRNf1s3zCF2TlGfRc0lMWmg1ymuApc25WyocpOWJQ8Gt3CWIUr7sfc
9sWSF8avvn3B/+oN68roLoibiCKCVDPKPmK1iHFMJfwt4Aw7dXyEIAJxCMsN3FiAtjPBuTTLbfUs
n0UcsXfmltNGIItZ9zunNguxyLnRnd/d5zwLd7mikmUHHpUYYh6MeOsHS1YsGM29plrHuWhMCIgq
jUaz97aexLnTdBppKL9yCkPKp7OQdws0KT5+VmobMV+ZkCn03v8pcYpgxrfTqlQfKNDdZ0kGazHG
qOZFcxBJ2rPKAGLMKAn73ARYm7eHmdxRf3EdYJkLcZ76kRi+QiX0LPulgZVeyy47+pSWzSxxAYXN
5LEDLly2yU8YNLvPDdVccySJqreG5WVkhkLENOKcFFzxa7zJq3dUCslZWTEbSuFr1NjNuRHDar+U
1eJLVqsyxrq/kkbjQGRydjs/4pFxVNynEKkuOdaaEtvV9yne4mVoYLIWVo4vwtBBvKcywl+soSUh
EWRwJysdVAAgAxZNuQUB6+PGNRFr6/PyBd8/ZSMlHeh+L3PFKc5Ao3VKT2eXrtxxoHKCp2Id/prD
pKZsLZWBw6zavsKcaIc6fEYdo0FiFymT67f1zegReyiwK1ZFJ2KwHbpsIE+HbfJZWYXIOh2OtBiY
O3BatjLc3fQgT4x1HlBeS2PbNrscvPjjhHaKjDOFJzODu3ZLhrpGlsHK6/9l93CJJ+XT3/y3mdJ1
o2Lbty37OjvsMK3liHdDsSUaCN3+JO+IYH3XfXBDOy1p65JAtFZuB2MMLfHo/aKYlJ/9c8uvNyTo
urq4ueb3v0wNKVI+pbR5P5EepV9HEPo/H4uy7cSPu5MXdIArZDBGQ8cupmhcRngvRLMqnRwDQOXN
B9FZTDJEr+JhAGRDt0hKNElBsc5q/UCHuDmbJbjr0d0EH+rz0odLTjYDye4KvV/xCtU/OJ7W5qwv
qXYwmy/hOLlInnOc9u5GZ5tY6+7tNce1cwzXgp30Z8ynjhWx2544y7G3UvyADGYtN7nMiuOMWsWb
kVYDxzbbMDDfXUlFPnTN/QhYmGA8o0rJ3tiiKPmRYtDvBhDr+3Bsk8o/f9PUTim5Us6FnDupHjBh
VKcO1TU4EJfIhIaKQrSCs1v0jawim8oLtJbjC+VES7DCrO5Q92RxqAeiqfsXVCr41KtmgisI6AKU
PNJUOodR0+RJvQRhL3NGwqROZatgkdZAKHhGWH6/j3xUnkayVGieXk9njduOF5WMYRWH9qlw3wNy
JQptGultrTlpR+27U12Y3iHDEWsyUABkHxsp4FXJsIURxuHeMjMjJX0fM9QDjq16jwK5Bjiy20Jj
x4lWCzCZgXDEhL/jJb6X3FmweVnHL6oKUR/PPNYcSaQSJ6Acs61F6BX+MoiwUkQ3cWiU+x06SPEm
Pwd9FHuBELOZ9aNoo48oFeDofLEIo/F7muhci5nl9xnRQjM5+y+Z/d5WFfZYW2s6qYfU8oUIgNyv
Da9mg6G44iYzF2JtJymzVa6beg+asAIYD9grqTFdS6XS7F6S24ft8cYnaYYXvnMiUzodjQOwhWxB
e0wterMaUTN/a2ON3iJJbsigEXkeEwLqL7iSud/rEWVFSJdVBA2Yvje/LnnuEm9FuW42vUauFCny
mmGQ/5v70EjOScMcmEI5AJ3Ajaph5oXe3gJ0MNP6fg9EfkdPS3imh20vRfDsMmTG5ga+dOpKy0gX
NM5lxCrwSPhctPRQdJo2sHkq2KtOwQ6tLbCym1GBUnmLiTcLhK2bX0oF09p3K56E73kQ2p6D8rOw
MIcY93WofsezFt7I7rNGzDkNpOR8srdWrg1oNLEtNyl3ExGmbboe2W/fTOZX2SeW58RMfvJ6DIrf
sVXY4vgrR/OdO3yTNKJrhYuZ/jG8nJ0fuyvd6udxIq+UP14Gis+KQ++Jac3E5EXgw3PVcCMSFIgS
OCL5sRFMAVKBGJHRo4NB6brBPQ+F9Ze2fwdMXB4WUt5hP0zAmCXB4BZGmgH3rwEuJmlGrCSQHKKk
jLRzBxJTm+3i6qCqRoxsqcvJc6EyvJeBQ0AjSNzjk2gldj18m7Yy7zH8fn9h30BMoKL1BHuKV3Ao
5NMZWGkO30sJq4HEgKQ09kKdfGa3iU/rUPxem7VYNxcimTJhkd/0ywh0y3FmhpGBsbuzW+2HDor/
C/Ar3Gey9ZxwIi2bt41itB8Y8/IkFVGjIqO9XBoRl7RvJkgdFMadmwChz5KRB2qRu92z1WJBREW+
q6M6dHn/wp+hShOfwIT5Wt9l/x/gKHdygLEAEGogV49KJBUqbjUAQwbuTt6JnQoM49JF14joafNr
/QSbgUz+BQ/aEciznymQ6xA/IjXhtQN4q0o4vyI/dUdlE0DraTmDILKdaDEjT8rqtEZCr/yXavGE
O16YNcsYdAFr5excvvC1NY02Kt5E8o4QJiGDL4NPAZIeB2ekkXb2jpsHME/AonNdXZRt1qiIF3ky
LL7nZmvDTPjgWem0JzErb2gG3VOkG5/ohfRhtPKrSFiHZlH1smFvYjCSly4NQwEcT1/F5DDEcxv1
7JgSXLzAYxPlzJ8WHhXJzt25Vt1/2eyqupukBmGS453fuHfr0RpGdjnDhLRggEoT+MFxP2bV6wN3
eyqnmm/I2m2KSKTVmaU3e+WvoLrFuX9WcCaPh7Y8ZIF0A8r4g4bt0ixhBkfzcIb2GPd9imuMyj2U
Cw/A2BFZOi7AzFtOJOwQpwVOl6BqBtzgyhcpo3DLiUWBzclmkL0oJTUauBZ90V60HZPPpJ2rIySr
H03DbiTd4YvvlKU0QYt6oG/fZcptC1qXemjViNEtmQa9RzHZU9RwuA39fFZwRUI1q7DHRXMnScYa
b1I8d6yBuuquLZbXSw+1z5xyBX7NHmvNFxwfufIIhYuNw04GtccwcgDET49qmNra26unY+CGFV78
yGo0rdLJwtfm5OlIyijcwzXXSivK2EjKnCaWljOcAM2LKyAmLwgJMda/gQYwh/EkkZOwwQwAsO5n
XQC1nO4b4+DpVUgyyPoSXNO6KSKRkLv1zogZEExHyPSIOY3VKN1xLH2nl6Aof1ZwTuZkMa+scVsh
trA2D3qyy8pePg5bQalvt3MPWPfj0Gum8XOe4HKU6iwrRLAmHOh4oD46RwVrBDAqbLDONay52rOP
plJdnxK4BSQyzJMDCuR8AW2AgY6c2lUUg/dqQPz7tKigMCcN49hGgb0O3WnzNJxoT3x2+n4yfwTM
BcBJWNb1yyBhTGRiJDTyC4NjcyJUVK+kgo4D3xcHMOa9D+j2EHaOFCvJA6bUjE6RLGhVpdiy/lC4
ly1tdVHMde6GEe3kOJY28goX0FiSgktHnfKfICoNA82MRjLs7KlEempg5JvsRlH5wRFrDGajGlWG
o3nWbLBlbR7Q4ssduN6AFi9107O8mphpCpFQJzDBJh984Wz4Kj1xrwQrKpPQXl2qPEKS9xYd3iX0
6/KjK8dF/XRX1GOywizD11bxHlG0AM/GKB5YsDa07t1dwe+RQGRf/k/OITD8UmefoqdVChNVrFcl
f1mE3HIUjA5m38Fg2bGh5BaiWfdoqgP9f4RmXQCvVMVmJvca6JConlhOgkuoeAtiRxJcL5IZk293
Q1QXgPo0GDMxLXDJD1D90AUIJMZWSJI8fqNhPpAxReHbKTsZ7xp21YCaEc3XB/PebOXGpJsIeStf
JTmcHfIGG+GQbhiwDy99PcnRLuqdiRFBMBeboJ8MAOYGD6bLQM55ftBtLtOmlZ9TDW9VBkrMjR+U
rkdiepz1fJ5wRBAE+Tz+AYbtMEJX+aB8KCSJIW7Fmz4IVF1+M4byn+9Wn7Dwv8C2kHjbSe/0pZIH
cyLtZgpk2mDosjkfi+BirPXYBx+NWW6lPdFSuefsDJF0tE3BIWCcBsEGZgomKM+H7TF1DMeoUNZn
8Byj6vvScPihWKfKQPFy0onfEu6WV1SLof1LzZ7qCXMn0uHnkSii5n+Yscusg+JzSoUQcJNk1JS1
XFlBPOcnH0FanA+YEa4b+6AANx+qTfodi2DHUOi4whA458HmRQTRXO7+RN6EVw5puuBMRE6zfeXp
FUAkh+q85Undkxfsbe5iPZcmO06HslC+df2TAZAKSaIjZ5k0l+4cyV31PYffjg8Qt8ZF5Ofm5F92
hTunJmBdTzDHZ07EGGK6wwngDRAZGPBXCft4+RG63BwaJquQEbwVyaTsyuUm3E4zlPvkQ3YkIR6q
aWzzvTIJcLkAoSsrGowlJ7LnioWvTpGtGGg4BZf+54YqJX5IW7/ZID5dddphfxA3ls3RXecUs0C/
2WKOKXaydgUnVTi7ltfHCGlj+emsKegjAU/rtesTEF5mHGJFa5OZLtA0RvPSf8i7OmlPdiyyCL9Q
AXizSZitWlSzb2E/n9E3x9v99ltT7BU91cMzRO8GJr8qW+ObO4OgajWTTG0rdGjsyJJcjZDkdeJ0
Zhb8GVmmC4ofyNUnMSLsyKqnBd9PxYukOznCmtzcSmdzceHHbpJlrnQbJ695TBkh2xo3UN1szGfc
DJBSTibKbxdgJ1zETbGJtQSHAlmf8jvv8BrTlTS5aSwKl6hNqCp70NeuZYJ5vj9fUFkGzEcKmQYc
ryT9ang7vyLmF+s/vmKXF1neKVcL81kBIDiwRKtalXnOjB7/eZnJJN9WccdbFiDCGCJTqct7fMvy
WXq2xuxxw2KSTh0nVTj8oRa1UnGcZTgn87JbQipp/dqpF6aS+SM4Qo/u2yiYmVNMdTu6qBIaaT/C
PDSIaq1NzHgu5Yvo6jZ8opzqsPhu9iegaonJlVJg1/8WC934vSVHwcaDCX63626R0JeNCWLsbD2H
KWPr50mjr/LWwfT5G3KV3OmRga5Pnf35CNPcgBKFHjA8bMSfN3r1NSn/lISGyjv6SV2Qr/kftNAu
PIzv5jzxUYLjLavlZ1kcF91uKgH/6uJXNrHf+aZq7qWMuhX6TWrUrFIDr7kx0/MhoR97Uv18ROkU
FIuHpBVXrRJD1Yoh+KTpeij2582S1/d500G0VOH9aa6gwqsr0sYyRxhFOnxvgZsBA2xR65lQPmhj
RU7e106AW1iCKiL+ZRP80r/QW2bDFCM7eR2B/A6LuXSqDxPuvhdP0z6XfXZwvzHLfBNjEmTJA2i2
6jSTPlJYjKfo88oXDA382ZxICCKcoN3/W6bK1RY8L1oDkTkAUn/hcdswQo2fgqBpXhjOTJRum8dy
PKihaUHG9EZOn6dlr6zocIlq5dMtEdx0qIdKK+7on0lCIrNsE5Yyt50q+L5WepnaPoj+wh+vO3w6
cCEhTUbvevPN/YFwsR/RkrZodDVWJU3N5WTTNAntOAIMgOiA5EEDWC1c7prxMAKOYk4GuUcgBKsa
BEu2snCJCdJiMOQP+zPrOZ9yr/1tEMvUfDDbfFfsXo6qI2D7nsZScrKlYFVFG8U/0XUe+jVXTEcZ
SDAJqrdW0mcVaKW1I8LRWTwgNvzd9S8W7SYLg3PsU+4rLZjIHwC9naIBCud2hEITU8hK+nqDfS+o
iWX7vjuPwCCLuVTMxFd5qtuMx01Fzxrz+FwM2lPGe4vSTMwKR3fWPbK7EinI0e8GKqi0CFAl0mR/
Qq0zF1UhpbnExUdaKmR9OHG0qTSI0zc/TFLU6VemtvSo2/uCK3EnhjSZ1ktjBfz1lzMhKzN1pfR1
BzZhqnZZ8B4RDsDUW3eiSiqfclG3tzrcMBF6yPiLfFR4gQjTGl6VfNmah9NzT1k2Zcvv42QJ3Vgu
l5A24auEtt5/uu9wL3yqAk5/jJPqHA295Xwkva9AKsfu2IT/I5Wt3kdiR07t8sjxY9hLNYBUUrk6
SdNX/BLxMHaj59Zhu39QEH3JAreb5UeMHxCR2Crqw9mBwcmTefSYwpvtoKpKxtTTT+ck1qS749vs
nXS9w/6vU1cEBh9AnaEszD1iQo2GBB2lQRTqzYwgZSw52pgTMz+z64DyO/g+vbUmfiqGqAe2Gqx/
+8+/89yzTGq6+TPY00GVVRr6MLQUPIX3ROkiipk/ANDchENIsN83cyRlfo7/yETD341uHuZaC/A4
pDq931g2M6XxHQqNstHjIyy2FppYaP6p77ltfRH12PcXT+RYlWfiGNteISzTprc+q2Lhaq3Mab85
1rh/b75U0OEB27m25AVxZF99On3wWkILBV+VJfnUARjxmMsiF96MBuVgJMrPvcH3WHIXLDO9zQN8
T/ByFTDmiLk089svxAIlgL687j/4xeJhbVq+mYBKZkbJbTEM0wxmF/SZCFkCr+DGz3s714uIFHqs
GABlee8vQ0pHR5mqquw+Om7YpmOZu1TsNCvpTtXstVD+q7LVxd+kH38MA3/ogtiEsofYuJyIRoa6
q5uxPXT3HcudJPB6hV0hYFXRgOv6ttZ5+ZLF8FvlnIBcA62uuiq8qEbE+OwSfSEdMCQgdHYZv+qV
SfjdkqUN188oiVcSmI/CMA3XxPhL9rpDNAyOOMOPEfBseIBnFJ2CeUf3ARRgeGqHGnMC8zWBMvUE
Y6M3+WUu6AQO9B4FlMu9S0Dr0wDKUK9JzoS75iIkJYUdvEATr+o7iKoXx6pPyKAQO1J+thLX7XLZ
bccL/nPnHWz0ZkbgnXuN9aBlZE0+3HvRMqVXnHJmPtogIr/e5ybqHiAFyYOLDos6xwkfwzA4wN0k
ZDLxx3s7eKobn9M1n5m8oTEsxV5Fnj6JOIzBpfekXWljlCaGw45MIsDkqJLHysv/4Z93Ugnz8gyt
UKwyWXarkeBdutk7euqN3noSm00S3YSpO75CGAaTASte7v/wZ561HMK7TIhgUyNQD6MJs05puGXY
us8h00ktfVcy1qGgGitLlDZaG3EtJ1aG03ONhoJxS4rrw0eqUM5Nupn/+KM0e0xpkXs0fV71YM57
1TwUFerecyDyHYcTvHozl0mwUxVpxpqSXy2stV4e5DuHbEJI2Wd1XXT1OcgNyWljJXUUeFum/WTQ
mHn7bVfiyrYX/sgTCNCblJtwp96/sPKrBLhvJIZaNXLw6Ib+2lZdT/GarsGUJM5KdsvRhxygM4Jk
FJVHyPLBtYavTNkBhUZjrxCgx1/+XjgDMIeoeC/n0R8EkjN6P/19WQdqmZk24GEx+jWvdSoTcia6
LlAt2a6H1hmxer9nRyzUeprkpm/Eh7w7RMpYLHuUbUWMkhrGaKx+kNbB/0hQxLs+RQxBhNqh51Xv
jv9MG53vuZf7bA2R/2KeL6Tay1R47xGrvQSN6lwvCPOt6SbYJfhMfdqtNR6TDXE1+7MpllEv0NHN
reSfvLSiL30LFMUIpfwzpQ24qMlF3SnZ9FlZl5z2oSgtNDnucN51/FY6MRVLrlztkjP18+JHD/wR
b9DZSxskT1FadlRJaq935Vq6rir5qfFjKvo3ufMgmd3IoPCTNQLKn5uXhfX2fpv9fog/PDxLzocs
bkMCKpy86J67BF6TQGjlq/F+2UjDHkitAsxUN0bzW5r8NhH3QAOeZGZZ2hIQAq8X6fper75/XVYq
+TTRpUwRSstu3Sx0BpuAm7rGB8b6KUZZ2b2gjSSbGUy12XKMfTgtL1JCOa5Is7hXjwB0gsR/wVYA
yzCi6nFm17JPQ52/TB2E8gx0YnNZbJKTCFH7Os9Dwdht1LAvvLxb9dm1bjImcl/V6rp096VAFQ+c
S2SbGpunriA6KM2/GzB37rr/ybMKSqPb7CfUC0C7yqroAIVZi3VIMVMsrE9ayfcSEThomZPvo7E1
VhyAuTG3HHzd6kbBvVC92XfTjgbdNiimuoiHdgFfdEUjswS/YFYDl41Ch+0VcyPMIdHq2isL56Pe
Xlmy5/r+88AZX0A+oNP2rdX9RNekt0OiBrxAly/DaKS282559Z39NbUa1oJlV9p3rAVuiir84XLa
MongSFhOq9eXGqQw7Nc4HYCVxN23Wib2nr19yDXKUDM45OocirWRtd//B0B7gbmqin5wFW5U0Xe1
DP6ylpa9qoFu93f/RmLlw3S7F2BbW30dL1jZC9rqoiynE2LJGQRiVcP76bpv4n91v1ZOj2IGpuOd
wlyWkUvHcMHePzUXtsmbyJuPV8wdW5SLQ6ypajXXsj6+xWlR2568S9yNbW3N+4ePT6DwKqML9FDN
Sr59VAbhaGTKD3iFyu2tW9CIvkbd1xc7uUZQ6AWSLetCqHVgnMWKwN+K47M7Mt6txqBnHNLn/0lb
/46JB8KihtiCdt3aCECqbmGED5yCLvGMrDUl6KZJz4hZ94OJYBzVjGtb/AFLKK3FJestlZXBP+3z
QGjg5ZW6ioYqxwl0OTYp6VIRK8fHkvMM6VeTaL/oftWAfTJAMbdVgvR9InUoiDnpk702XVNomZ/f
zWpb9kkdpqWqjcaJBx5heKVvBcSDeLGhthBKZnANimyBUis8PRgh9hHOR9+W9+IP7RgEn+IWjDlc
1+MsrkJGXhKNajkw3cLDKNW5gQwRbvDEHKGmeZvnB6DQICRCfMYqZ1n01mfOJVI8Pii3LJHsAEP4
SxlnZ2u/OBVpCD2MQER4fm2hx+i5WMV39okmaGQgHrh6LQz2tRjDUQ5HE+bY5yVC3/qlJyQs3zQd
mZLkIZItL+ZnFmGchmwggxoVNTJCs1hG6+Ps1G24zPVoPbUW7FFslhV16YCeFvYRtx/UtoPjIajB
W/a9b2f0R04mErnSVah6M+ef/JSnED0RfNGO6vPBjPyihipeE6L/Slo8r/vlFu7G94g1IthveG9u
6By+b+HkJy9YjNIMDINnBqELSTimt6DX2HxwauoYdkM9WDD7xkZ3EMUqXIF9ar0Dgx4UI8FZSKID
DvNJL/m+MK3ZmXEBEruWRmM845ViHWlcxJP6MJTgIQRZ/CX/uEUuyxqzB8vY/03vbANJB9Sa2D9V
lSyDqqUShWc6eUwser4sgA5tVijLnhLQw170zphBanokwHFXpcd3Wh/9I7BJAwlq9ICR38i4gTkW
JzqOl9DlAfpTyXTNp4V8edJuAoSG7YcykwzHVb6ZrdCdJoU5YNNOV+IF/biyMkvYv1Vht+dChoX/
zVL4M9aNwDLJlox+JUtO7Mi5NyMR+x4FgIYVRSLb8mLvuNR5Z55erhAd/BM607MZuiqrC79ZVeRY
TP8879lcnEH06Kd0Ow4K7HDjh4dNyamVIt4+zHAt+Yp/XWprcjFDlsNkMqsxnF33wJUoZoXgxpO5
Ke7t5lkhwSLiNUVR8X6p8AfyCF1uV3XyMMdu00XzaDy45YrC0We8dSoI3+w+XANvmSMg00CNX6Yg
VKHFQCTc7C0rLf7NFe9cMUgJFBSbHWkLGN4SASvN3vaYSLiLn2VgsjxVj5+TXkr8zB6sDCyIcznV
yYQc3Q2dFHnDdHhhJKIo9+5Y10PXKFPiiFf5lHHKlz8Igv2XtYqiBqeKmBuwMvuVKSTHZs6qveGt
Z3tRUuSDviOjcLlDv2kdi8PSRqoucp+YTTGL2vmRNlANkEYXDQn+vyIDem/DmPkDGCMPMQu1Nxqg
N4t0DbvBZm4YVTUuN2k+QSL05G9t5S+pcyJuhzZRORdqLapr5pSfDBC1pGXXcF0FewxdQHwa7AZ+
vyl+6bVMJ1i0XjzHiuPpHar6ajqVwgIhyV8x1GbH/z6lS0nlCW5VRHz2g9FR5Fl0flHVN9CDoMJJ
PRgVEP6wAHy+qJJq/XvdRg++zo/mik18YfincNaJ9KXJ1iZ7bQKazhx3F4lIMq9D0qqpXIaC6WwO
v6VeaQGPZ4CMRYsELYEg3Pjt/Y9B6aPjFTnXpBKE9Z9z31yw3o5xBetnmuBohU9A3ywPGe3kbgHw
ESfx+LW4mdAGqKKA5i/eFdRj8u5pgneIPvomGD3PQBkWqw9687LmpBD+hb4Dn8IL/UllmoThPrg6
HpHnnbPaXbDUuyCIzYgTUiEF4Fwjh8m/1jP1S0rVHUCwOLjVXpRLTIJp1RHYeBcABVVi1eappges
d2mCNDdrNdupf2dblX8sSnY5ze1pVp+JhV/N5jb/UGHxIm0ajUiLVqM6KFgGRpyxqSDUr8eqXUcv
eOmrazexEap9+ccV4iO77NPBrRJBnc2nrnmL1ZU4S40pznKSY7qHtXcaPDWcmmo56hFCsPpwy8uQ
GCnyIjYwvC0atIv+g0URmKe/X0fIxfRzdT51wMGH6KHxvruomqN9A7B08NEnu6Epm+bm7kphJIt8
LWcaoDmpI35FfsKfJA8H37ExNMxtUma/lceprflZNMGpPpHdPO2I72T9YyBD1asfZCy/X5lN8AXL
40nCzz+W5bYm9tHAXXDUldDH7klxek5EBXomUAgoubQU246FHlG0ijK0UMcVhv2f6PRyFe1GsTDA
+SBnnlHDd64iMNWAqtoX3MIEJey3R8hDw19vDHsDS8jaUlIOv/Mz1MU7n5/AvcqB8Guf2mnrZLLY
i+Y85yBzojd8IIE5VYSYVUiQN7jlRxDL0eQtM7CHh5AhP5tuXOhUVRTxfeG1YmtWWt+JytTvla8c
fXwI2AqpyBhhzeZopl16xCuJqoGoMUC3vTfP/N+xMCVJPVCRJq6/5FVwqHXuiUOTfwV0acWUXa3F
SeVSRDz3fO+h+2ixKLgMFiFpaoex200LyW7RMlKXsAst87x6EatEHoHU2wbcoMkLRpo3rs6fVKbx
Z2sIUBatrqEFNKSA1QLFJSOej8ZDoPHJWZya9PwEzF8VRxVW1kO2fQ3GQ8cAT4ZxvqTZo/CqX7tt
pOHqfP2O9Bc5Zk1k3tgkYAIs86PpBAW7j/LlJaRz1opVOWVfSMfsqaasbDgpkxJmBqAQ3GH6+Lab
pMDOJ9Bf8JOSrXDxeej53r03Vix8vAMFO/18zYfS6RRqy/KfzhRZBfJYhn/G6j4vu3yG5E9rFeTK
nwmX1cXUiLvHeYApniyuvMJGSoxXSZ1uMk5Oi9oRP1f+qB8XIaBeJWyl6FWoewFY2sIqzidJ4DQL
yZ7hmvA5uT12T7vVANyJntKC7QwIOCMfIH4N20yprLtny/Nq6sVAnuVfUTRIlJ/YUoZr4sq0LYRs
kFWwSzPmeWin7Ia1sKGb3D7RSjN/cWe4YXgjZI+MnA0INcX/MJNw7dmFSHWR7ssPtdMQUuenQlvO
BViVV6B5aTxIHVVHFthzEezJQd3/o1PpKw8iGBq9DFVRrr9Rk6YxyyrsCO2GVCWhaoaQh2kicqaB
1mf7tWZQvHUMYa85nJ34pga7EVah4AzcG6oqsoC5tcjPOpMXwvASOjvbQq3kWPVs44ejS2GF6yPZ
HjHzonrc3tesaPhiBTftz36OMNEgDs9zJjNK1W5CW/g+7j1iQWQAiQKahrtUgIuWqSvvpAJVFRYM
eK7HUXH+fYF0jLi5ppQB/Huns9XdihMNC2N7P7MANtWIoEaW2wevRS9A0yWx+16j7OrtWh64CFs2
2EEzQVaIQth7LOYKWO6aurKOsOGfO0IagjvnS6OW3Jq1DMGUwRkfBGQfSWfOVU0rjCN8YIQrPvmi
j8gaONO1Zn58ET8i5mBOt5qHfQbBV2JgNaTiAejnpQFJlD048eRyKEwOEyYuV7V/U16/TbLWqU84
+1RX1CxzPHc7T6g4ZK0O27CupxFqDE/MD30QLh/sz8rcnSbQYKBS+2/vF31GA3cKi1Z5IzGx4t56
0VYKDj8rSt2HLGfT5OA5TE5Xwhn0jtMTtb3CW3aIruemwriPGSfeESarQooAdn2/DBmYsOJZ4G6v
6oX6qBUTY6JSmdkRBCSKtg4xnRwpQyOKweI8rAFOSpS6GPmjtsT483b2+pqxP1g11KTxR9yXeiis
M6gmL3x7r9iwZabPEI7jYLjvcwoVB4chDosGZE1cWlsbOiHYxYqMx7UtOA6h37bI1k6EfJvwvyid
5Kvzf33ZLeDbBS2ESAR+4/rj8neDNyP68zDW1acg8XFhJIqab1b7G3YhKaf18wT4xIcr6n3JLhQ2
/WugDy/dmqE9wko1256hNJ7mBuJNv4JfBwZlz+0ABqGi4A6KsosohDFMqPeve71ssdB0pB70MBIX
5t5JVTa4Y4O7rRymVcv4wt1paJCQDVHi+BZfCYigQrCMjWzj8BUZRiqv8v4wxlpQXvdU+3ok4IFC
6BaPaxH87M3NzvraIMIZ0PLxIhRM2HuzDneBymv33t6upcXKI+EkSUu5CyD4iGoofcsqtSsPx3bU
GJYki5heyNhQayg1UoLbxy67JCoR2V4GaHy4xRSvZZsIm4bNRY8S/nzeV56AJOowd2Sa5tEoUbc2
lN6THJYZQ1zStntgCI6eYSX9im5SOMwMpTBDLrsEr6nFKOkUMv7IJqAxbBk31cGrjrhr5/Bm9XYX
iD9iDxsNbqPgUPMmAGSjPCXYt+ynh26TXI13roGEcyCV3CNBUaO3+xotu6CqSWTk/P8vnGA1gt7o
dzIELzdl+1Sv5DIzGj+YGJq6rvDalJeHuDc16cJTTR8aGPRJKRxHhOMUL2IavBBA0OF9COycoiom
EceBD+yLdBkKhZ0dxSPwZlSNiAI/0WLEwbN8RE4Mqe453y1HAChEcCLSTnXq9POvD1VdLyFOmXcX
SIMbJWoiS+ZqpLGK8uI5mz9HQQMIFzJQjo5SouNCv2yz1LDvFej8iIRpp+YOQqVLMa8zwW3T2U0h
jgNxtWQSqn5ghxpusOu63MP7h4YHrdu4uD+/fqEETOHOgFYy1/okjp1bkOklxVjpMfR+7VsTXTDK
nvO2vFKepguLbJMRBy0JVDXfbC0D/PxldmC2fkCzo8cQtCk7hQvYntMEoJCg26tlEmx6/JnYKRAU
w4fmxomMN8oFrYlwA03Q+iR5a3PaphiyYW81wRwgei3qe/AUvK0+XPVIOQM/rN/F+qEx/Ajj6Wb5
Q4bpsQjBqvqcgVxoB3EQQdpmwwIfm1lngZRWv5p3ei0n54YSdvlYKhcQS336sryyTKtBLWgXFJHp
OloQzmcAvcYrg8hYZDAjGqcsAlKCE7FQPqk3tB3D2IspYv7add78JLh6X++uGtlGS4FbKAuJCir7
VCSIxxjR6CydTbEXtyOkqYvkhJeCJWYi1p2Wbg+pai0K4EcI5y2I3RA2MVAl4S2ZS5jfAvxDvY+Z
at8nOqg9KQs4cTSwxlobRX7fzdLqcxePouPtYa4GqkTzvnkSzRLdph9jZbMztCx6FEwg8dCQ8PLh
DQ+SHPTqVMJ3UEvz7bWJ9ERrOXpn+eC45QdjPli35FYrEZ7BhfkJg4E6KjVDTtHas3aRunVBxmA4
giGFV02ap0vEJeNTco7dSlIvYB5Eq4uf+UDMzBNkLVbiJx+gwJUSNPsPco371x1J9PNd/0+a2KH1
GGsEXxdyO29XBgHy1N+v1gUyzsxR1AsKaESqQl57W1Hm213P9GClGBTjsmGrlE59QzEE/NQ9bJG7
AlIM0gs5n43bOwCYYStK8p5GkbF41rutismai4wKzIm1yKtHiZSxquSEmBhCkYvgBdXutJiv1iZG
FZ5nB0qASmM43CGp339K14ZWJUZhX0I/RivpBM7HjWO7AriDEvYZMh0OnJc1bfnG1m5dLo2As3FU
Y8Iv5Y60Z4EsD6a+bCWPh1xWTq3EuZMlSXEYrc3GZzEa6ghULlrWicxNZ+EGVUuNatQ+jkWjNuYx
drUfRsl61K/nJZGvOKQPkmTtgZl90nIIHLsAcri5DL5rgViFPpQAY9mBXnGwWDyMJQ+yTVh/Vu/5
VdSOUiIfedbMufa7LduG72JfIDsZn01eW/e3FICX4du2Nz8cmoeiEi7N0hW8F0Kk/Hn3rKE6W4i5
8bhBd1FpH4V3S0P7nhofmdBgxqvlKdT7XibN5H+4/CLW4DcwDSJ6QovN99HhIEOUDlkxwf0rlHE9
Qrp0phFRGzvF4iX4weZa5L4xn5/sBTEP9DeY0U44xjp0zGIKoDrvko6j4vVPtJKvTCDB0fQ6D7Ov
uLgECuRN6ZY0Viq4hA7NnVE9MaUc236L97G6Ab7YKuO/yygDVRV4XuoqJHxb2YsNZIIv8EAVbmHT
hO5+zQrfcKA+K4/IGojd3Kc28M9CfxOHnfxbw5WXbu0EmgruMtka1hOuLqXSyZhYHLbywmYttQOo
W1ZSPRFa2hMdFwpmaqKK7MrjUTf/ckh1oJhiuzvm6PEd4tHdq1WriqyV0mHoD1Ss6QKQCohJu0vM
NxNXhXi+0YCnaMihlYsHym/WX2JXxk7zxu0tZH423kuva2rE2sG/nFiPc0FyT/1A5E8fuOObQ7Va
SGpYBpnQdsrumGvGmJg+QRLPoQBCH7MjbC89qZciNnsX6mVVk9fCu2HpaD78ElVdRNNfpkob4m7k
jS5OX2D6X6VpY/HioBHejo+VSrz8AIqK/7DmSHucO2thXybCyWk0HPW7cpcK2rnXW01l3xNC0T6m
J+BnqO6xLHqixDGd2fsdyJbfHDmZtQseCvAezuJlvVSvQ7z9yF72NwDH5NcRvM1usCch7FpoXgkc
JCxsZLBOaUl7Pgw5UcGZKh12QrS9uIOHihdRY8ghOap+segV7S62kCqEWg5F8Mzfl8xrvkHdXYos
AKV1vx3gEaJxRFeKNq63HzaTl8wWYX4uTOQJ70Iuy6KxFKBtjONdzHQRmzFjuhYQWSPygMqx6636
E6YuSBilH7484hcIhTg2rdZg/YpzaXbSnC6wVtkH9Lx2FwGAAU6uFc+26bU05QMCsbCM5i98ZF/k
QtOkPXrPBFd07aLcPy3X+uS5p9ztDJa4oAiq/plI+n/a04jf2wIUiag9QW0otGyJkS3STZN0g1uJ
pdxvYLg/s1eNnGrbtk4ypdCPWECKdl0wwmP/y0YbjXfGF4pPAO7w/L9nFIUxsmT8v/evrRw6ff/3
BQIM7XXp8JuvAHTP5m9pv+ZoGsC4dKDAWDtlaCtkPL+Ir8PXCQZw0IwrVuVZjQBAE1fr0hAa+ohn
T3giiz5enyXtz75HjRuUUTrisey2lx3INIr6QKnxDeAFO8266I3C2Tcx2tkXSN2xh5V/1HC9/hP1
XCtVQK8JmSw79Ijim/vAqmg4aZoImiro/QcYnrDO3fz6bFIMR0dYV9MfJQwYhsS/ve0aoylHNay4
ew/TBOluJ3uTJ0Vi79AG62rEryNa/jzUFLnPzowUDCwqyZsBndfNYmsL/9Z8mvUa8VTLq37lNSZd
8+SwV1ZS7otfeCaLNRbwqsPdxHxsobIRzCg2/zZLHZJWV86CEfhJx5vZ38IyEHha0S3ld9uZ1dkn
wKmwuidmQM0sJoVRMTj/9EY/+y7Ndfy4x0b+cexRjPWGiHx66tmlUYGumKfeeKuruIdyVSk7F8PT
2fZbpuNqXZVvO0Vfi4MvLdwkw4bDg2ao2yNkckIwMxfk66E5s4sa+5a+0RfA2xeO10de1XzOS4bp
VfG2q4Q4iVSUlwOba6XOVuucMqEHShLKcGDjCWAnD1iRvPiwn070pUL7K2PVZ96fc/puh8NUJ66T
4wKGuajxlMe9CM+Rapchf7guh07belujyqhKx7u+wWMDansC570JzyhfliIu24fIJU4VgoSw94rq
E3u0I/AKkHqNvIMXv/vk/SYij/PBH6at22xnIOwaN88v0g+WBS32HmgdAzZKPind8bjk/8Twe3s7
hLTlnmj0JG/fSlVqwDn1MBUvCC2OYelD0KvG67nniKDcKHUUVt/PZEXOtvSXhTn5th/MquZB4zC3
qrKHO4IGxdYMKxtwZ+4vd76e+nuMbErb3Hh2kbvkOssLNBXnUL8CI1RhIGhG+rYyW4IrW9CN4ZD1
tcfvHBiA/ZyPoS99+w2gouKprVzdIdK1wFQzWTynU7DVieeHGY7iHDyE21eDE5TUde1tY15KN6Oe
PILhetGuKoTi7HnTdKxmY/TOhv4KXQCkolwVDH3H0SC7THRohyx9RmL3GRvsW6UwEknVV14S6lTs
9YWqAER5aFkZu0y/Er3kz6nuSXVWTqX95FDV/39+u0C/soxmj3CZoPOqlCyWZVItKDm9b+P8PKuU
w5g6SaML3hYnwzjCo2M+zYxmw+1dqovl+t8qk+/HsZ5a9dESuecNJo/Bz5vFmPv0vewugUW6kO/t
DfYfvyHkO48Kcm4/LWx7HUPUye3rjAja8jA/rZgdD/kFybR/WgzON/8ybnQRIU3BSqrDSMSPfkbP
UFLQy7N2199ssXs/3GMTKMiXzsXavXXQYtk9xwqCyr3Xy0h7U2kF78aT1edzd9VA4zLCdF9LIIb5
Bzd315d4cAfJVWRoeRqqm7P45F8iQ5v0ndLT/mm4U9V4HswAd33b5A45fUwD6Sz243NnvnOcQvH1
CC5jIPgaogVsTeMCd21H861vALcHJ76GvVQdVR2BIAQvL1dwPk7mDb6j0i28ttkk7Bi5leNDZC2g
rEUdRmY5dPfTZgPiJGFkteNFcgbYDP7nLuxfBX6tpI7rNrlnW9FKKP/MfU6kuO6KMeOANHegTbbX
3embdw2nhXi4R6He+xtr+HK2HEoOgasv0cZkecJp2Mshe87TZK6mM6RvdEgKC9r7AleZeiPcXWAj
sn6+gomjEyPsF71AZTFrc4QwmNmAxJHLvQYadKhqwZlcOQabslXRATJ/Y4P1udRo83ogBfK0uDaN
tcgPPPhc2Ymmc3fSIczmHZanMIObUUKGggcabf9JwplUX7MTDnzYHeEnO05DUq1u8uTZF0CvNeDz
jqh304/zmnam8FUpwAwy6eoU6x1KOK/Wm3Gh2oGiAon548dxOD5pHi7wDVVLcveO9jGqdaXfg4Zl
++/ue/8FZxpleuUSobvqsypaotOichu4K/5OyCnn2h+lOZrr1Um1piGYni/Rd71MELaS2oXy1Np+
/dOzhXY2Os0F8ITFyFFRfast5vlsiEp3QVhPTxUE1gzYgzGDHIdDFlYoN9AfP3qpixJ8Gi90CbwT
QlK2zrPuFswZTUqR5l+ALli9hxJMtThe1fIhXhCTQWW9It8qLDY+JfqBXBefxwUrQJZK4qqN5XhJ
Q1N1YgBsQfFm/j+C+exOem1UTC5AyR3tQWlZxJzvWRTmbR72zybJUZ0OtOzbDIzEeRKvdArj0UKx
axzPH03NVBbH0sRxzJXYe3O9JN9z2H+zQ6NREoCYSpESWV9TnVlNGYD3hBjA648cA+UPtQORiJsj
CFLC6BqzaDDHoar5xfEo+5v6Gq7OXgOyZS3YFkWqKNyTfpnofYfAzV9NEYpTJIH1hWAHqoiF7Cuf
6Odbt4I3Fq+JlpZiMzm03K3+3PD2kOy4RdtwIOlA5agPuXYzKjzQhKOWipphD1jB/V40N8SUbA6+
rSfDbt8pPE2/UTcP7uTZuhjXjCjUHRhjG1nGBoBP9r/sddyXl1kxPQMlnPYy0A8RpH48P20egUX4
4sMIigJ97DHbzc4HTf/yhY3Oc6KsPuWFSNUw4+jMr+8OhZX2zZPnD2UzJxLjmpIQZ//lz0ZeF76z
pvu1dFTDVT2b9reja4jAh3rMY1yyY6LcTcuatnATtIehp8i1puAiXFbm5SUp+Wqr6WoUc4fafuB4
1LuWsClTV+dUGLG/u8FBb6Ief9vuh1PiluzRiU/QkUkvvnT4bbY/5MCa6ye7FSQUl6bYVMWRmuL7
4jAOKwvHOf2jY8EjlynTa8HUBPxS5z4QopBmXNk1q3Ma7EATPOfbPasftYATgh0s7JHRHwX5Jj4t
WwQ2CcgSjS0sMtAXt1VpgGdZYxw6IZDtYHgCkdYqTHdOsA8LfK6tKcYKxK2JI61rsscMh//B4LCQ
PABKn5eGDNrQG2xsmBTPW/cMy60/iH5bhkGNVQUpi008p2MyiRffrxwCa7+A0wmAp2q2pV0n9sVN
6VeqbYukb06tjLL+mC3ibYajSt2X603SsBpEpv2Igqshprwpm3IqYyBAUiLOGp3ZBFX1f9IoOAzf
N+HxuhO3I1rxAwzt9ZHz6IHOTrj0kgEIb0+n9225XeG8wfMVmzWGgX2eTnHz1sjxH98vI82hj7uz
0dIgYgKJpAVCTLIB9d5UQId3qTY7Nsw33HBEBAUkn7+IJW0nKnpM9723DISekSET1/vIV3kwsBCk
b4eNm7gAykr2qRSDo686jpUNPIJrgMQddoSI3hKSs8qrJX6BgjccljOP0N8j/ok1ZWIEec4edOQx
GRS2YGfVAPU2U2HLrhcy6wwOpuv9JwZqjvGloepJ3N5iEcw/qRT5iB05Q2RboWMuvq38PqkfmF8X
yb9v7Qh2ot7Ii2+0U5iSip+xzMkNt+nErC8G+yP1j/UjtcCA/ERvmC5XdLMpM286EkY5rHQQ7QmQ
aVyYAFlck05I0NpWFbleoVt6di5r7hKo30IFB6/hpxMoMRWxdU4aGx/lxPF11+oryd3ajXr1eIrq
zvTfUrnPztPmdbLpICqrwYa7w3/5ObYpW+B2U2c4hB2mIeNgNJTXnRzhrPJNVLCONRkoiQdel9ge
lDkiW0kR3yv9WL18ngpuWRqSlWsWbhmc8p7hPivxBBaJhbBMj5fORwRnZ9QmQDikdGI/IaWjaDgi
JmuRNpLyd6TA8bd9T3G975Ixbzd2wXzG6zFYRNlJBTpUPOrAlgHW0T7E1h6H5IqnHigBX1SmxPvN
rXsklQK2NjDxzEscSbnz2Ca4UwdK0N0MFyt/gKKn+pMXRXjgKhlERBkCqbTVg6HpSuwQ0pvdMbnC
RAyTZvIdVvo9CSNEHNIctELpXRDI509JRo9x2DS5Hjezpcr+Kt1cxIP8cKKiWo0cxq9jnXfHuKnQ
mot9CUhHw8uKVWva0cVdwOLALOe+Ze4pQU82ErSsqrofzKX7XQQN39304mHQnGY5til2TYnaUr2L
+gXAJ/mtZ/95l/bPTSA4OpsPgHTWHZBnAdmjC9SFXssI65ll8xzk/uRy+jIiT10PSS+Pi+3JSVWB
7qjwbQYeaTfn+I9frzgJTjrYP5Dmd6CHnokDBnDNX4j4u+RT2FtmxSWLWDgjp49nxTCf/dF9wa1m
SeDwT4mpHS8foUppOVAbQ+8Sy0VzTzZFbpPgIktJuB4rExlCvNCZCSiL/Gv0I5W+kUVcb1+LVKAL
I8ffxr//RzrioY0UnhQuDsnVuX1iHzcPQL1K6kUYAY13kIDsohQyqFwJnmqZV7cswsJ8S7CHYa7e
cpD+2o5KSyz1EeWIKc2+31kHEFCpImxHvwqXncJ7BnoVRpq2vY7T0nSZJAxp6ueor3HQtvYpWd0d
Dor5NC4H0SMWK11eD071NP9BflWHIAC8Um4LLM2gEU0KUyIy08I2IO4F18jJEvjNg+Mpc4ryyrt5
Pc0N3gtA48uCUPJkcDV+mT4qWiI1bL7CwQGjWwy211qauNIQnR70otpiOhPfuIY1Ca6Q+6hTTNVh
zKfkbI+R0RSzDJXpSEPyf6mM3T55gue32oaSLqBn6ToOvTlw78n4gOCHTZxHipvZv/K4OJGR0Yms
AqMDUfuttoVJMu6QNBFmMo2zmbwRYDJSeXet9jC8ie6Wm0bYyK/75JUzsVlBFT+YTrtUA2jy8mbN
+tLbtYH6jau9MfJHv1Gu8cPW1WWPysmVouitZW1umKxYgdWQ5sd2VTkeJKf5NZXORKnlTPPHklP3
3xm2meB2POybMsim1w3bz8AOFD9k5bY0EeSHs/7UlNS5FE3sjOi0+Z3seMucDN8ublmtlrcC1WKC
NwU6Pcb1/RWkU4smyfRStdfZuvj9EC+rJ+LpUuBJ/1HsbuWV54oUPq0ys3wwZE3D0npdofXqVHq6
b0T30g/dqDEETXMNKYF/yJlA0JqB6R0pwJaqGSJUblq0qgW1bcQAN2z1h2ZqTQ5UBt78Os9pKyVK
/DNg7URqfnUd73tls05JisurP0CM5pIUNlJi0bohEI12epPmfKocaApKdI849lLwNmh2iN83LQti
1g6mTmyy3cHJHHCJJ0+j0xRnwCXagX1Tn7GKuNReSOUsnwsMJLZEXRoq2c1XdCmqn2a32dMqjYha
hDSzhfv2hqgun8NDrKl4BW1BlVDRFp0f7d3ME2kGujO+Zr73RiPHlc3jlzetCgg6rXxHtU9E1m98
wtujw2CITJ9e9nNN1EkxY7tO8X8wCGoCR5HG2Zn2W7K7QRr2HrUkkjPwmcRj/VgHN3ZYwWz2w56D
vwGsbACrKXQEe1ORhf0x+gMMTf2f3JWXV/RM1WdfKl1nhBOVFZakKtLf1dJpEqZujdWlgya1NYYI
mhVTXqenBjVFY39aczbLs7Q2u2dL4/bqUzb1pLoqvQXGW1cOVkEDebToSNZq0XL57B1mNYP8h0nL
ZCFLSxTJD6aOgWlbm0NKOHys+z1Mm7m9zlxHr5U5MRB8eCnFjlAPa/La0j9XIjZDymzFcCPmuiSu
P5QDIDUqrKk/jrbtWxAo0F8CCD9xEOTaCLkZ28P9tSfuExrBIhxxTqmwTq1ep9Re0eKDGeg/PCPm
Ns4Ds/BMZ7wSyOzCxIDExLqSmo8u5LJ/c3wMuT9lut5TcysJIdMVBtUPFEUIQCBjbq/B9S/Z1c1y
NnmU2+0WSFY3BO8Befo4L2Wu7UL/EPEuqSfC/N01MbxTwhGSzy/ytGN5GYrFA1MQDcTbSTuWt8xY
RbtO3bX4QWvn4mgUNdv1Fv+1KNVdnSXrWS1gPdBf0EvXWidMo/xtoRCZoV6GPFEkYB6OBdze5SFr
bdKbxYVfBb16CCy7cjTRuxr6ymAl7VSyLuCaMpjJF6unddICkRI+2czH/hybQbcXgzbw+PWKDHIV
zDACvNYIRXzyPeJLiEVWeYHmKmdf5QTo4VPNFK3sXZeayFBZPqHZrFrcxuk1z7yMw4EiJHuR5ZKH
ZxkroqFw1kXpkg0fNQnR5T2RfNzv8uC8a5zaKcKq0yW1t2qJa5mV43LokNxuYeQz7NeAwFmqBdcw
lTUT31hDyasdRO3Oj77rXVNu8sivKDK8wcjSmwu3ptdGlibCsUghNMJf4BzOgyG+uXJ4H2vkh8ko
Pa4iAASV2ATyJQ4LUStZ5GXtc8sLXLb+8UJ/lKVvEaNYNOm9YxO7ZonC8dwXyqeOnzNpr4IgdAvS
PCqBnKD75utebSjkf0hpk5T0NvZK1jfwLYdM+Rav6OQy2QLBIgB1s31Iv8FtyTxc3LHt+q9i6G5G
Sfc7ljH0mtQpijc8OpAN4jiItmGLy/n2VncveMXDZUlzwTp5I19lLBn99SmudjP7629nFFitYxA1
nkZnZD0ThAXVADlHLUJQ5nJK2iMvWNe4zQ8QHkrnRnisDYNJ9HyxTsUKKKayrmI6f4QUhMs9/BZP
CuITiGtJd+0D9uJfqxJrkcdjcW5tiiJ6J08K49wJjlOraErq47jti9vrIEu53j2v7EXXztgKSvqS
zcKSmugZiLZ2b7jzAZQgAIg3E6Bn3Qf7l7TOgqneNzBDA6xnWok/g/BmnOpmfzhTI7bJixMvZGdQ
oAhmt5nWDc7eIUi3GuakofEUwiWXcTrFbq97KZQLuxCrpIOABd9QhqKHLJZkdXdswpeFUDv6E6N7
4WebPhXgf7kwDExLNBi6bQffljO3fDB+9mjS8cUfbGWJTdH4nxRf3Z1cHod5gB4LLFFooocyCnVy
1SesZBBel0Z1yCDrVJbV4otaH+IbzNyzAwJQB9N/eCiqBQJ+2LGJpXOUAJqmXHPFL75kEnUtWp2b
VPsX0RkZhXKgP3neWf6MRZrMWt0fIBeh324J6g5Y9Uvu50E1zfGl+HlzIy9P19a0yARTSOh9a1Ob
m6fiPmpJMZW+3xcojDk7k4bgx9ClO4QLI1E1bOL4YE8RG+WcyIqpIQptktSS+SHpB9UKPXOyYcXM
RYu7srbSWAeE3aRnQFyZEY9Ny9YcxUECeLKWVO6iODzWzvyeia+4IcVppm1Ud1fWGOIX+Br65kpb
ACl+3P2l8tTex7HEgb0O0BHY1ULEp6vdAlhkqhHzaIqcx7JaS3L0vRDd8VzB0V2wqjLfMxAPEMoo
GXhxGzi9sP/B43rgn4zM0VPl+OqlEFCGjQGUOqNIq6gDhU+LaO+BRoURCiVCvyWrJW+GPcGxuQq/
qk3fLYac+yn7AZb2uyvgId+7JkwT9uwRmYOIsxOxs6by9Ja31Qt2ZAYWpXrpX/kIDcvyp6PDfwSo
naonQ+GGD/NU2XGXSdsqO1e/1Dlt/3PhYaHOb2DXkSKibGY8lvrtpZTmby3LsEKxwZEk/BkXjARa
3i1IoH4bXKikwCQvl+DDuN+n2Sqn9czyW0Nk6gz0rQiB9/V58Diuj8jvHuuxICsAyG+5KnbVmNC/
kjA0/y0HzYvrL3rWBfSw5Uv3uRI3i5W668v6JnKzfVx29TKTsj3hwOoWBulIjA2h0XXGhcOfesKU
wr9/mpqv6AOuQR/ypWzh9mUyJ0i+IbTBRWmWZsbI2UXNpavXWfWn+5820zrrs+TwVQdGnh6x/oa4
kDjJoqw2aGYeucfXIM+toxDj0PvJVjGSs1rpTIk/Po5CT/1ckmQqpNN2imWrDVbmXvX1L8rJ0CNk
BuUNRA/glDw1vXXGefEH/jSiJ3kY2qyZ27Bxz9ynP5RpiPoxMBcLv2DKRimASS4l7e6LUFL61cOZ
CFQxXOg3fSaE7BoXcFnZI8Y5hiswWGFgswEPuf7HB5lribERH6HUVL8clJ25Yfrf6AcNVNtzjjIw
XiKsc0pugvYL3EPP6k0+tYgc9PHXMS7qfFyMgB8fFIgcoHeWhuN6evVW5v8cHTVsqahyzoyeb29v
3bWRwH6OOwRy2LqyOe7+X2+aTloQVyGTwga7z0kTw+XfSXG86YwaAp32wmfnkH6B2esbs1UbOGDC
xJ4Xz/UB6Ze43yc4TjCPh+KwRg+ynwrZbmyNpEqtP4zQaVNV1+b8RsataYZjBcpFWVx3AVMICzPh
ZD0GPS6r1PiUB00RuxeB07wXdYviazcwo3RzlrF8WCQOWlcEa5OBi++kc3KeQe4vGFz4MaRag82W
MRlM/LV0MUKYvmCZ4RWX2SpXZ9P7Oh5bgByYy/qfLeI5eO8djmO6oCI0vYT8MS3U25hLg4DaPVEQ
N+w7IAu0gTgPv9rWIEaZIw4faPVIv7SqDqANhvL7Pu5w1GXppnLZlppzOBDPioxMUbLy9HSXJnCT
0lck1WP5HJwC0NtUhx3QrJZyNbajZXRG5/k2TLl2CL0vt9HX7ioQPUp9+91xMDJL1TNHzuAjTlUS
waK9+FnBaCzWknny86CgsRNuycNyNQyOt54VvukZ6HLfqozdXiKB0cze/+y/FAy6ujGKQEYxsIxQ
Oz/MzinCnCUXzodxq5PPKKRSbJb1WOxEASamVajnOCtDod9oGj7XjNkuxz04cdE+dxJhq5Fc5oVQ
qdAyJfZPtUarqngFsuF6NEwcytD9gZoY67oLpynot5N4uLZ07iYj7N5IrfHmDSscjpyiBPoTJCo7
Hoy5VjxEnho5f6WXmUUgG6LRPx/KRljoU/bqFcRGwZzjJNWsZKarmsNKBiKo9503bkM+fVY91S47
hLP4sKQAG3Uc2mNMBXfvGi9qXQOQh6oLshRY1Lx5+vfX36mdpW6rnVgAoEnppDBP5yzjwuY3YZw8
eXLXVj556VAktN+OxDPi1UZao2D0Tw3/8/eTt2Y0CUi5H20jZjYknnpQFk/BQ09iNnvry7Xagljq
uxxDnQqYieMS8qFSFDRgDNuRua6tOfFtP/fEEAEb84N8YPKNoONFXBIC28WvvtGwtBpDZ5NDOH/4
8rJQIZYGDnFRKjEDE5V6CPjIvbUA1lVUzwpbYOdLyiXAJBSfJz1Hdi0RooOyht5rn3UC7i+QuUnE
VWsxuE3aieBjxJodpXaWHngj4Fbq1WojBhQmWDQsrtv5g6RoqYBoG9d++HIjK0s5cGajfNr9KM1A
VuWdj7yK/3SMT4XjI9u/r7DnWBHdo5zU0RcKxvkIy6JDrd+7+erae5FgbdL+9GA0f2y96k+UBXi0
MFjS14Devy0vRYX+SLtv/ofgSGSvE6r4NiPKreWHczNEvB1Q+THouZFraFSYp4g9RraE/QhVo5uc
++/TdrO639J8nEePTXZeg9zHMScLOnDcoHK37hHb84IG25DmyvtTo/nVdYU5qe/FotSPLui5b/8N
y7bkr8afiakcceHp867ZXFwJ3/iRVx/T3GhmwMNPDJRB/AfOzuGAbC7BkKks8eMLfu0XB9MYSns8
1Djk2Pwd3WsFUpWaWhy0+sFjoXZSV/XLUoc+RaOPiJU0k9DVBAkeAQa0bF9M2BOhVKF75Xhkn/ME
0ManmdfdDe4GPY70FLYdczF9v99YdMtbMQXtGcRgo9YIJ8gyBxHXIOK5GvWkRwDvAhDTvf1HIesk
arySdxV3YASE2i/ZDOxdCcUHkJFQVJFIT2u7t9hvyUD5CxsUIX/4RgaVK9HIhiAq/yNOq3yYlCcS
fqjeMYomBlG+1aQ7BQH4UBCdR9U1ysPVKM+muvSHdJ2q/sN48UophnjkUDwERvxiQzDIahgFz58b
s/SZyeH4WTaW5uTvR95ENX2DLrY34hBOUg8plgExcrRP9uwywiVKBEpJZzmS+soMmfWEuFPZKhxm
fSSI6YK1beEwwDUfY8FP4/IbKClYDwIEiRvJ4ofpQsfH6PYoTMxjSmADnVPF0san+x7ZRQQpcOp0
dNMpDMQntlOZtoQzyn/QHhZkdSpyBwCAGQYPWPKxpfq8g49tL54xlnKLzw3NKhiaAVlLzDx3o10U
F5kObpLFa2a9u7G5u9x6DsW/s9R0iAiH7kiyr8QaEGOdNzzbf9tmjEFmY1TI+2HsxLPa2SX7ZMlT
8JdA9ivfvw6j6j6qC4ECO2i4CGgo7VB2aYQ5JNoSKMSPBDSeDcyEbPryenQ3igYpEZbNQq0IBFs/
o5oyjGb9HVNpNk8SPz2t4QPxJzo2vJnPvmtv+GiCdMwE+RLbetJTR4bWH/JhsrB7oHJh8EROv9hr
PxuvIY0pVn/luAC6uwOwbO7DZGiNUkxAud2wNj51031q8+64NLh1F9q0cO5V9HUPCtha93oObMPG
KvURWKSsWHX4D1q49Sr0lalRG7EvOurtz+J927kMIysimFd1elEjxwU2zLIEUnRuliJDTQpLwpDs
X0K1foYEkiNpgmk/VctAJmTB6Fp6GQoUxEUhQBkHUZ38gBfvqoiYnh/qIld+pdI95z5i6UHh0eSp
C0hBcpIQa8VlGlZHe7HiOwECRYirCXKHs74KaulFZm+0R8DEo+0793SuxzyYfvdy6F2a2PnDgv0F
4fOYyYBKpqIz6sqnOthodSWHk+eopWlqPsK7bDnC3SyAHtMQCx534i5yemQdxgXohb2/5E8fv7UJ
9EGRf6/huIKFbAf91RBzmppRfWofi/JZ36q5n/3Gw+gjc9v+3zQ48AOkJNHzwyIzq37ZQDfhcby4
AUTZYi5arLc7NRk2ayNLZKRL46gyveXJL3w+8PCfEPHzJ1ayzdWiIB8SEXLD7na+Wiq8/FnzHz3E
DyYtaAXuha3ucI3FvgysFRFiZLSVhRTbykwRhuXqB2q13or9XLDiBdNQAswIxP38PPrU6mQ85Tgz
pD3UI5ROvCP9BTmgAUFUWTQCBuh6gZXYTlZCD0HVQ+DmiTWcfw/ccMeQqv1m0nuTClUuhKoNHdoe
oKsJAbIiAM/0hdtC3M0HktebSSgyALiPakA3t2+cD6OD00ar3EckZ7+elAmtRNFcyADL2OsQh5qN
Fw1lUQUEyrLl2ORHzBVtR3tmkkTv7gC/NutTkVq2E7H0RI+qYg2qcQnGsySjoty5sNyqQ+fASP+Z
LNG4NmD0PQCQgNhuMXJ5fLmDdBxX5PHpKY8FUipPKuiohMWqfPki0YOut3szU0jIx9YAsN350GEh
e2xYV+SU8uQrVzHEf73BIbcMVf3chYYpfCwUiVL6sfXS9hCSVWIpwZd5k9VAaqp5o1opy/tTNAzD
jMY4SLPnMhOQ+Q/T255jp8IHdz5hJjkKomVLlFXm8CA3HXuOxlN6SxlMY8FMb0S6u3UMjn6sphVi
cQxukOb7CC7G7WeIzncRabyaLwVM87IXQSppyD5KhTBwhebmumi0lnICvySzJkm4kSjt7rhXH8QS
CFKERAvA5Was8cHBJsNMHgAwXSF4Rlf3CQwxLufbw54cyz7qhUHJIbVWpx/Y3LSlVwJgixNHWpNN
ntSpS0u9KKBpwxVFgRlfxvz90m/e7R3+dRe9T9JLrULMnlQBJO2IRT14yK20Xu5U5QEcZzYveGKh
XF+mQ+M8ViuPkUr9QanOGd7bteufSGNY7B8lcBnPf2g1fYFiWQfZxaT/A7GHb50YpM7xA5cbggUK
FGef4FD8oV1EmRPa9Nd1ZuVCOZUAg/fNKX1+dccadd9rB4QfoiqnIld5yj6CsfM/yiiGkKY36YPU
Prroe+qwb61Y/RuNBi5XDkI9+xQ14xnjYihba1sSLWPMJv26Nhb3J47N7N4azHz3keHc4Xd/OcWb
tV08bUbtfQP9mnj0DbbHxE+ZugZqZnH0TZlp72IZ8InepY1oAZFHoTbLjlZU1ITi0mxnixETTY6O
Cxusw9W4KIjvdMm/G8C9dJhSFpm94PXWzfXpcjbluYxtgB06eFUslWrRmM0OLEMZS616XWpFoWQf
sLYZnnrAGMvq1W/yKBUD/sce3K4Z7LPRhrzYrpsxseFl0TqVmRdq0K8JWBkAuGt1iB4DRglVbwpk
UJO3TaKnn65ka1rFmVCp8xeumEX2srU2pqdxjI4CYoiSn9F7mVu+29VtUyQy39joRKoMz0lCdjSx
IjYzw7WwNpfbXFziB45xcnmGscZ6eiytDpLMVhjGb0hdQQEDidf4R3WGFzIAXn6UQXe8jtvmeTg8
yQfwjkPlDZIgjCPLFvz0wNoocZE7dr0QJhYLlntEi5/7ASX5S2Q4TX8YgeRx9fWF3A75AFKNu+h4
nWwkD70PKNs837gFe5OfwY67Jd82S8gZDBtLdxkKVj8u0RWQAbxoKMKRfTSPtf4ac8pR2DmBGdXd
cZSI/b5JQKaPrClnFnYHQLvRvohKVreJQeR7y2tBiGWwelmXVWYdcginEWt9dZpJ8hS+HaVoxKTK
o2ad56650CjV0mz8bW/5rD2ODbH3IRw2AN7EZ2akPYz8ksP9H5uUSK5Mc5sqcS25t/5Am7D27Tj5
7Qz/HQzX7UQhRY5HHvggcR86uuBIXy8Kjkcoz4DhKfFgbEBNG8+XRv0n0rFzkQZoOfeWq0XbBkil
2gs8aVpykpNnr3sLVrnAuDQegHT3p8EGiSrjSVzNzOF3RM1f2O84Bzr1F4WZbcTNnG+Oyrq6WWVT
HMuZa4KIavmPilkXqdVlfpGX20yX1YJAn7svhKcF3bClSD0FMQeJMKH53OgqgNQOjR3utABdfxn1
biBjx0WL7pdbhhipzF233fDWXI/TbBNWjOg9gI72x6K1X8nBU0P+NbFINnmWRLLgezu2nGKIEKcy
095gEnWOj4J0qanqhFUl5tKsQybYou26cq+KVObRP/xCoclkpX7Zb0QMUx2/v8SqU+PERoWHZeUc
9qzeU464/Xx4gIuiWQPXrbkEqm/6KUAEjodyiY9kCa+XfgLoMfzt+2UkSa/l16JK+LnkIklOoQio
Kz+peBbgJnlw6pyQ3Ql8xhQi5ZGXM2pX2V9ZgwEYxWra9A39Wnj5wWPIhp6D9MVbtS/XuHI1cyBJ
VPvVTADIZaUIkplQyFC0mVKbKfi91CdXkydCCFr51EDdQdlHDhjg/bqsSc6JD0BJCQOH8pxsw8jx
GSiEUQOa26H3DVqR66gmoETLNHsbrw8GcUiYzFiI6lsRdQWKaImkNuBxkVRpAnyst0sN9G/Xe2zD
UwMGdTG+KeciKe93cQXcXreroEwgrsmqFXd+MmAmmTSZohLvDNqrWL4TG81C65LmFIgGaxxDXVsV
RquVRkNqE6+eaw7P0pWnzVWmB3lbj76g2d1sqcLv6TCylxVRy/p4+zNeRRBTL6JMz0eW4dJTE9pS
cpJwSJqGcn9ZljZ2OaQftE21SBHoTcUVOnrr+0mJ61NT22nNiZdLJldfduyfWKrlM0G+zeNgxJIs
MyccYvTVda7jC/QnJXii2xbchRViE/Xko04Cht9XkIh1vKerSg0WVuWGHwYeOb06I+UJTnQ4CWmb
Paypgf5vyzuSUFEZseuJLQILT0j7XTEqGy3Cu+2ECqDW8mSi8o1ENDEDhfCUu2Gap2F8gJJtd8NN
zfPcSfLxGAB5ynp/Lf8kyiX/PVfMJI5FfsmCPn40NSyRZH4er6XXU8lRF6q94waRfQ0nWDaHmS+V
Dfb20HFARApdKVl0UVKzGwcLNCOVmyTlcdfiJ/n36pp7ZtEhqdKcH8acuxbnB/4PZa/i7wtaPRgr
6cmv8EtLGfnUiglnb5ouyIIkkDNUfAO7Q5dMjWQynrWGGyGin8/nsbp3ilDgtcMpSNpVu8O5jABM
SjUeksUnjIn4jZxBoHvqggZZd7eR2p0jlTPLHiC3fLXAko6OE15EqQsNtGivi2TxGY1PCAvXuWse
JiakKX9x7r/lUyLAEDen6/s9Sb/3pJBS7hCBNh50qSh+YGnXIWo6Wu8xnYP/OgkIKByBDMPUKKaQ
MjQA/J7G/3s0FyTFFXrzj1jh+vLJvhGfR4yYE+McNliqiNnj47jqDTWMS0keMVfTTEuXXWbYFsnB
+bVN1x5FiYI3lYgtXsi1DNcR/L3fBNJMVJrNOtHVtDKTKEdB4KhqJAv1nnEIq4hL8WJZy68Dmxlf
0Ys8kJ1DIoGyDtyxEok6M4cW2KiChipnX2cJ5sTS46yB4M4XFp5I1dPU4iH98FIiiAouCA/lBE1K
7IEON6EUDBf9cBANDgWyL2qDRs44i6b9J3c5+yQt0SNpCvdYbw17wRNw1L0UiEDvXFagQ6mqL5lj
spxRP1AeFxEFYv8GcfF6rCkXqzTQu/Gbxtwe34xa86dElcXvQISIHyA6Kno762OAoCL0Pv8qJ5kH
QWRAI5nsfD5PV1o9Dh+GAr0phIP8u5M82NBvvZQeCioqht0yUVeXTOSLtSqkZjeyCnxSIj10DKvA
rkROSzg4dVXruXF57V2AeUPqp8V01MR7uiNwujSXekoxKIjtC7FP+fjzspYbjUt4HDbxRAztzDXK
DZDrAmgLSBa4ywa+l1IoeZu64Wt0l76YKfL4AKTdhojd4MK8DlBYusM4tuiJmNhh8OAMDmyUN1lN
mcVTH7qJzWdNoH/a3phdn5JPq+go5Ton7NqbPzBmce31EKAoYi2ewvgdjTbjFdIiaxAUblNjV7Vm
UIn5bwKiwcT0mgYpjrIqrxGWGeKNJrefcsN52tetJsD1BaC1Srz3KQSj44FZYpPQseZE1cP7n0/P
Li5y6kYR3CYHvTu10397CucTVg8pXK+OX5J8a5QVF7/LmKv2OYuRNwvBkGX/dmA2fwf56/HPp4Lm
9Vul7Tmd1iqSDEz666nW7fkMMuBkGu4l89nudZx40/a714jf/TPV/brx1jrFnFUoStJK7yKfuYXg
PXunJLYS//6ONupptuT0tUx+FYRRUz9z292Z4s5m5jVJgwReaJ+uECBMHukzw8ONFYhBdYb2R3X/
7uQHwFKL7nLEFGbY5KNKhjyvO36zJ2HfD8g1DEc0TdX5D9ia0UWipUcZNXegs79VkeTniYj8aATv
FTR+2uh/p2EkDMXjFpJc4OZRsXbZBYmykfbI9vOkPMJBVWfiY/lZwg25cEmCui8dg+XYKR/ed9R0
Miu47OQUvRQw8EwdsXyLO/HpPM3KmEJsKvz5BIDxJ3actGXiVdAWLgHDU4sON+0Msfdj3phC0h5g
Yk4BsFkpzFoAWVwGfzgDqGuX/HPGD0O3tI8SnsJnsvp2rJrc+9gAK/o7lAFl+gMXTi6o8ywuNxk1
WaycO8t9AwevYzTGvE612QB1NXmaWZy3Q62uTuTUyDjWdiMiy140xpwbaRob+4dpuvX2rnNOhPCI
QSZM/XJ1b6oElXACne51UIxRG71Lw8EGKovn2AxEzgY6oA35/z99DJ/mc9mVZXTAyq6xi2+w/iRr
uNSlwKl85qHnKF3PNYFM7KV/hnLg8T4R1wsjpDCjjCidLU3x/xgw5X966hO6Ur/J6MZ09FY3nv6z
CIL628FWQcdchOvQ4ZN1BXD4C+PiMIJ1MnFArUsa4iusY+z+BfdnB1/OHVXavvdzk9fU+hFiQHSp
d9YB5M4fTaBIbrgkbd2rZuUDlPEsAeFaQSq0PKHUE1k/xriu2hMOlgreMgZMCNkmskiaItF8GAfL
e5TMY3Kr78gRQ1+AuLbTXHsJe7PLXFArWiEM8DFASdPr8tRwcri1xn6TqU+PHP3MDZ/5yrPs0Nq3
c3g38vm/CHijjN7yoz06MvUz+2v5iK3vtnwugkFQy5IAaoCMcpQ3p3ziSI0kGzAnpDOjBUeh1Pnn
t077n+Eg8con08OjwYPfh00AuZIXX5u5eyxtIl1CjPl6aYHeHGC05j4UrbU+kjNWc7e/PVqL7Gbh
8pn11k0FuS/tumrX59EkzWpsBfseik5j9x9OQiWcolImF6mTTPUn235FUvrXBUUUS2nk6oYW4Z++
p3zTss4wExeFLcNlahKaLVEC6GLFB1pcXw5OUtUKLj0zjsgW4JuS+ka3oPXJwJ+kDrbvItonwleR
oUTuZjchT9rGmIZSA9TEyE8a2YPGqbzPbpZiECWZwktRaYycsngmoxEl3NSGGQJzD+/eflDlKv+R
C6zhP4CaYvRU4wAWYNDvym5+/6q9uo1xa+cG2eS4bRSh5DGtrXk2WyNHsXObrAgpZxeLv/2j5l9R
gEnUrDZaG6KFpZs1uNBSf8krefMad6XiF/QLeeTvi61NXSSJcDqqcU6kWm0Zrjf745uJ52VyG6tT
vsBDlgjC0Cj5fU/Mhc7OdYWYuvmzxUATidLbo7/wgw605V6v7lnzvbN5gOJ9lYL/EY9cytHQ4XFR
ztRuo5UJaVwVbSjWVGt5C3DVZDEDZYX/AihVpscSujlKb++ZOeDOmWQP+DRcNJCjb135cvc6L4Nx
VI9/pMJz+IThoCsSyKWZSjmwklzzjbUKkksGMXfvYfAA0UWzcNrIdv/DSspUWaXtUSnW8X9HjG3n
74DWCftpK9nxauhOQujdDZpxaOUXHGJdyWx13XAih8A5zsQ1hZFyO4PfXvwXOGExTO4eH8jq8U4M
Soth79GS8B8a3yS/jBl0CIqjFzcb0F8fkKFBjv6uGqqLP2Y+2pgzzJksaFkcy5WXXbz8O6B2RMPb
p7/vj/Gfhvr1AUUO2GfPRv9cqfaao3xrUHKsudXokgLASKStb7eCnOiSzuIbWyL75x+MJ0VFl7fk
JrXItoaq0hKNpoNzeEelnr3KUcpH59U4VdEDaEFa/kGHg5GIxCcRYsCLFWnN+t3eF0AQpkzKLNRK
jEX09tE7FMNctZG0mboKRr1IqlTfWb3PNk2Gcb9AUFwYSgK9QbBuHIqdEkFF+A22UjD95elkxIae
D4dcmCFnRtfYK0Mh/AyYGZZucwCIHivpLv6IoqEHk0ksyP11BwdFbky9DXQlFdBu+A17zz76x572
4cxOhTk/r3rhd8ls8x1IlmNrINa11fBcXDi09Yr5s4gpePodt/vUdsl6PKUe8HPBT225DDEPSwol
G/Q1VkQ9uoYc5Z8rHkIO2hzn/qmVQkmxbHrwXO2/rg53J332nT4TlIazK7kEaaRf91yhM8YRfyAB
pQZcvVWPpRk7+fDKxM4w3XLOK2eFwApp3QMATt195fVoPGtWVdJ7Txo+K2Nq2EobfYYdvO1+A/BJ
MVGS1psSs10VcwtzKKQFPt/Z1Aq58id4TwXGMamFuW7+laMuWyLOoqmMbLTY/hh5xn8rxfjXMfq0
CjRmw220gVCWLqrRuTBW/oXhlaFyXLjSVDhfuUFuy03wDlGMGEqlZwi68NxI+kfSKaULJHmB1hxo
02FxF9OZp2oWg9hm+LwFloh9LjpefIcb7gYUAD5H+07rYHMK3C8QoeOj+hyf7atfW+ocFee3qVkw
AO4IdJ4lebq/mSOJT03dMjScsGjM0G7ml5AutsTMZKowMDqUTCF2JVcScLFftvHFFHryAQv5onh6
GOj9c/szSDa/jryPyww8gwPmm3DZZlqVhusp2cLIrZKY6VU/LVlx0BP2wVGuy1DAyBy3VPRrjFhV
G9cfCu2v6tGYXsVBLglLINNtcTcB41WrkP+5dFUKi74XsJuuCqkvrNhVT9kQGGDbz85B2+eUUBNL
9pYCG58hoDvMU1orafbCpsDQ1RX02ELrfq6WGkWNGorq4Y4ruCkdk1IaFgNcsfX3M+gi2T6GFMV3
+gmo+e/ouErwcCXdWf3zz2fQFg0ZsRq1iFd8GtWjXdq2nB+Qb+gT06IaF+/cdEEebchK6N1QOk5Z
9rxDPy8z2Npk5PVVgz99wzsaUfGOO2V04NChbKsxGLd2lJB58fm986smotoML67rtaDn5/PkSMXx
+eIA+Q1ldWWRuoR1r+U4GXcmLxVzGTH8P1bdOK5KE8ftOTzzNxp6rMnUlAZMXAn4bB/22fr6NNPk
qUOVyA20QXqQvdNq1hjLlSDbBxBZX0oPsPrXPhi0DbcRGPbYjT0RDX4doMk0wMjJermV0F55viqy
dVb7jpKapnzaHbWeZAHwM50kYxhERAhupvDoWVGLHZwnpA3IsxoNu5HkrEkVFd+TTWxUXSEvW4Qm
XshZcaRMUMjNQajKZo8wEEDkjwpAuehlJ53IrUMU3xieR9ZvTpAM8WMGh92HC/+WtqGeEOT5bsV0
+4F/HT3KwIlB76MgBBAq7kbizEttFO2EjAkq66sWwY1LDn4EDhFIpKxHbPVk+my94wnzF1wELsb2
SXNF0dg9pG9LfvlUAWEsYPb9EOXQeLrbmI1Yp80Ik6WaMOnl30sDhsSud9auPrq5YABNFqpo8ZSu
+T6+KaRvTnFnwMZ1VQuVXyC+lV3jTM/cBmRS5HDLvRlZXzuLK5A6plqSN3OeopzuKPiM0x1wW8pW
LZZy7mXlqyImbuwcgFsl3/GwX8CT0H1GEeblfA1A7sFstdpZL13x42JuD5KAFcQD6prx8DeDdJCV
c1giL3uR256eKSEO64sjpjrUvnIRg/ODbmVAQv7Jt3DmGRC8xD805k2Sw8Ay0QZwNWT7fzgDB2aA
Epoa2clTojmoCNNXvF7x1BPP66XYJlrMkjmfrbJjxPtNeSe4CEVtoG+4foAYmdawZlT6TSSGGB2Q
RY3Nf0nE1qVfZq9USiRkSlJNSu1Ts+acCuXR898qbMaC5teAoprkajT8RkfaTz2ePDw6r75GBOBQ
td80drWehulmBL21emxDMhaA3zly/zYnLaCrPUo74j0xIDWRJS+QOe675SKMB553VuqXZmhR3CtD
n1f94HEZ86x65tRYNPbuF9fAu9RM6UEwYgZmKDb7sPzrZrNLl1nt5GHfn2N/biCZ/BOrNCDl7YRy
ipYlEshpwAigDIetv13Je32H/uG1MRFzkPIe4sQ5+nwXy1Rx3Rk1Xu0YuFoG6hH1niBrV1LyBPKr
PHTOYw0B8cakKaRRRJ6+VsKJPreTBNjv9Zvr0X2jkzoalKG4n3oKGlOmEZgnU9svvFd1FvTdJ9Jg
PeDhXpZkgrycIQjBoExAzIK+6nnLoTisuGzRPPiTtFa1Ppq8J2wVCR/ASlUC2zAlVU2SkKUAqKYJ
aTreLJIHu8/42wxg1W1042IqBm43aVRSJioBO6QewsDBLbKCzGRxn0GxtK6QY4i+iUIxkuesJWvY
QB591t0+m5/3A4YrUgWMaN6iJ4T7QZonxwmpcBN8waKFN/SXdGZ7Qa7LrWYS9/GpSmwBtuxEaq77
/wjCFtORXWlfYrhOAN3gQiTQ29qb3K0RF/9Ppf90TgUc34J7F8Iw40F36l7H5w4wy1ESWPbREYa7
lyCNlZom6UL2ej76z8teMp8plAPF5QZSs3eIR2SmMaI9iKR+6T63JPGdtfLvCdhaNXY5FZk6JaJc
hHGbU10CxpDL//CJOuqFDNunBkNLgg4V3ocyJDTTjeAvqSVrslFzbXXbRY+zuw0Bu9I2U0LclTRk
yH2akg492ZBFu3Mc6usDnap0k2YtgXahHEfOygSFTMNZufKkh5vR25W59ldBAntCQi4C2NjPmUjE
LG3KPXwg9a0O+5w0j1hOR2x5RLSt7Ds+RVi6v21LCgCE1JswzGbJ3Ymg6YilvD5NYkIhR2JFahYU
n1kI34/Z83f4qIouINQVs6hPndw2W4k81jMDzn761O77qLnRAoC7JX0g8a6il1FxpS7Zw7NVPxNQ
VKbvRq5wlzxKRKGsI5H3Qa/1XGq6Lc0ytoc/S2yurvGcFVwOzip37QaIAfilWzpiDFtEzL0xrLAo
MeUYed7ZMzSH26lcpXkKRnnKAPxXZHNFwGf5ikq/8CDMZB4rKn+gHeY6Rdu2fTg/IsFmiT7Dtimm
ewMy3ONRunZgCiXuWe4ewHTA/R1GpvN1AyELLh0TzuvxGIP3/UB/zwR6ScBocHjKNLrBGkyadTIY
7NDtnyy/saq6LgGKMJiPoviVYwx6zYD2Xef1qLTAH5iP8Ro2jXH1QYVZYf4eaQXV2gW0tC38XEbQ
mJBxbnixyUKtVVgUmq/gAuR5Gtj9Nsz0VBGSpM+2T36KNREDkCmD/VgxbZoP44g+PWze/cPCT66K
HtUNleFKk7EO/rY8eyVYRXEUEllaLxfvHNkbM1tb7qNaQjynXrOvlTbUr/mPP43XeVmJrNIjkM/U
7i4bHuawGkIj8BzbCLKcqWfUKAKwl5rrBe1Q5L75iwpvoI2YzK/HpEJ/skRxTW6eLWMCs68CMJ2D
qi6YHDh2IB98JHuEDvRUmNb5cibFAZ7M8xXqrJWjyt8kmaK0lnOtkTmEQqys9Cs83z6W8G3q+5zm
EZA+5gblOqGn+O4pHrfvZ649JK/f157UMUeMTJELgySiJHnU2CEBu60uaGsc2PRJFyR4oH0fo1H+
pz/SMR2ZbhtR+Q3lO+72I5XgRRV1ts+MG4ypMh8n8IE3r+H9E/Wqj4iUdRmdXIwKklpfCBh7vN13
ELkVwz77X9P9rsg5Sf9pSkdACdZ1ywoKZQHGTJKbxJWMQ0lgAO/yClpoKQmF9e/jIcQjwfg84hhA
POdRJKPJrDKqDdB2dTyBTlXMIQBU84orL11RRoxGvzsPIAGQMxbzMEwjq6buyqW0w7X+7P/Ar146
RIYrVruCE/J0Gz3whr9fvFDF/wjwYNo4fbiWLBqlMewdZgLfpTs3grv/hmjrn6VeB1DCoGKIWQyv
IGZQXXCK6LqiNlH+qLQIQvR1nTg+GlqrzUA4vWOs4Wua6jv6NsLk032djEs8+7F46FsGQERcqaq4
Tl+96ct3e99RNlLVuZ9dD8ym784KiIf9aF/7iK88g/KEt0SFtLBoVVZMIt3ytGGEq9/0y5HOn4Fi
iWSnRcMkhDPdwkXKR642eE0VZ+LtW/IG8512bshQ3XdiYuvRF3A0505bxVSRlGRUV+mY1l6dq78O
KQAk8WJkkiKKOss4aWMrVNKlIxF/5sAzr0qGVAwYnwpKxWPDUAn+58DPcPR8bft5Ge0obRoMq/jW
/2Rm0Rw5K+eoP4iPEDmhAtEZ/kGHO3LISleslQCL5oCCt3WSzokMmxEriu+v6qDupCiazjrf1jZH
6f8AIFjJCbulHrzLW4GlbfAlQL4i4jjYNKOjKonqMlTd+Du3HyoM9w33eHx3rVExYg6JUapRrcfP
8RYwR2QbEZDif4isTYqN0UR9cwKdxxGn4reNOOmJYcla/1/zgD4q/k0V2SFNEZj9ZAGjN+O/tfxK
TPXAd3mg0FC8Avm9cSk8+KIwBAoWPGX++HG3PNM+LNAzO37k65d7GINp3ZRQTo5IbQg+a+EKtzoV
LqS9L3FbMeF625Z1cAawV17Ue4UNNOYwh2mX40YiLf1hCGhkd7SESzgldSZ/40ibv+QGJ0I7sya2
/uBkPJw2Qama20jOdg7ebvcDykcPZ65IPDrFKrvkhNGFRVC+C6r5csVC43ZC3I/lBb0l0gQD7mIt
3LJ7y8F8Lw50hWUGenfOq16+bUldcmU2ip2y2mcRj6pfGotVN4kfCcqKiAHTD/bMCz7+F/WwA1/6
dpAsDlF2kFK10FDVseLUCKoFspu+0Ufs8cxxCPBrz+NmzVfteEUaFjakPGeFuoKZaRYG2fmk7cfr
ikGa5jgLYvpcodLG6uWHkc2HL3WeVcUNUeR3+2rmhG0b2n59kVrJqdBGFYEyB+aHqtIPBVi9cw7A
9ZVCW+PXER6diPyk8FB+JCwuhb7Nk0+/Qgi54i47cp8ydVqzW+pTs//MJUUmeJLdRfdL1mEeFERp
04jfw2/SVjQTt6nOFfsBzeUBH/pyn4WJCqmW+/XT9byLdx23AYGrgtBqv100Ajt768XqsgUXImdn
jTuazeWIACQaP0u2pAzgxkL+h5PJJoooy5FvCoufBGmkiUnF7IUluzS4bSdCEVcJHFE2OEeUHxt1
56riJEmmOXyhk45tLJjNxf13fnEgQaZ8F/JCQLKhUvyc0B8nLwlXvDMdzh+glFRHEVCc0ow79HUm
CBuiIwjxK1Lkw5kzfvCgsgd2ahIWcQf/i0mldW5VkBltoYZ/N6WA3A1J0B0ANj+vQbo66EbInv2c
PDmAS0IE+5DQP9YzXK5AiOrTcKYSC0uy9xp0reLnUZHyrJhwT/wWnXpK/v4jAJR7u6YmWK/ytR1r
kpu4K7QJQm5HrOWqTsX7ASSphwXqtgmip04XtyxJwUPqw0+RKBWHXUTvJUHjbROdDMJYxWNjNoWg
Lh19gZtSq1CjXdXjn6zhOyfknuIrJqh32TaeCQx4wHMQqQ6Hh3ZpSiOpR3t9xZdNAQeNoBsar6cx
rSNpalQH4MXrNezbEg1Po4Zs1+GEbaE4leW8A7lxRmnLuJnLyTZbI8cccHsiRE5pFIEvfKZF6BVj
dzX9tFxbLBhNcFU6+LD1oaIg8ZRlfutXMMuQa7q5uG+oRbNnYwH8ZTQJFJJ6u0DagRqDv+4d3ccS
KIWrHOvUfp5oR6wKD9etk/YcgXepxS4eWFqUzyjORveVCia+b+1DJSdsMD4mu6PdNXad42wIRpHV
4SgDoPvmHBDv91WI8VWya12bos81sur9cSxKu+LhI2YL+xp7Bp1WbO7yeU73yNKmpqF2Fpco/H7W
BOa10ouC+UNmEbtWkeZ/RZqNobldFaeICyi5O3dmwlr0Ey6L9QnC1GqL2/y5YdlIX5y182Rwtj6g
KBYJunL66W8w7wnB5G3QRUNNdX9yR+Q0TdYT8zbpVY8IwDEvMpyNHQg208h81ndXaFBJU9qxKeZJ
pp1N4glRFkHgjrcJIhzlt4joHRk3A/RYegY8RcQuwQaaPwOIPwnwYeDhwfqRLwS5v9UZRePHyz79
Hz/JWdhhraId9mfn8vHgDKu+nGTMnx7817V/TwRqmabnYW99IkXKTxpOSftvKFaLkztZEw8ftIpV
Po01hOOQsC7JMqOugyw7q/IFME1hhYThgDMu87vMBm5K1pJy41yN7L7jrfWXTCke9ZAQytVaZedS
+JNqzNu2a29szy1/8/xSuiT4neTbhctWcoQdb+zfQ9OiR9JDjPPvgLhG1B4br0uL5vQTAg0s4hgP
CyiAQQgFq9NIIntrgP3EbDAnfJJwqUm8KCRrKq2M75D81+6qE+EmoRG/rr/A8TyYjwfffq7EZJ9l
XSG/lvZsxqODs2DoAJ9qpdH3wITsU+JaB36g4NtvFoEyHLxYRdvzLKOfLGoF0nxO8aw75sEtB4Q7
SMkHiOf4SPhXktesbQCC7Lh7Vz2A3R8J7EnzuAx4W1VCg6ZXI3SmqnHDmpc4a55TE7ysWn4QEYwA
zbEygYcsQXXIr+MARbgOWcGSnuYGgU8quPPPPJV7bk2+/tEpJP2Qqw5Ub3zYRlijwZUmwOZDgVw0
2+Tzd7xdGhfAbn29629CYCO9owy+WSBbgnkp795CRij9T1/fjaM+Hd9TKRYqMwx3AXtoPbH90qRZ
7uzeWOo1IEcY3kohLwjSxQinqAb+tg+4uW5jTe7aD/jJXq/YY9Y1HKhdoq8izXc9FTFnufQjVIkF
pUQIJFr7Ikev2WuATwieLnmzgkad/xhlpoPAUepsadEeOpDzLj8Ca2i4l2ZRQFQLumcPHCxYcJje
PHUt9St2Hv4fFDb+LuZVz+7c3pthyT/R5v0wOnB65EAYHEkulpWz66D/laxPiesjKPQ1PYw26ZHb
ghe82BhriReAnpyW3UpmChQW00GlyflABRjTlTfL3voFeNevcO3/DWEdfFTe3NBs4X0Aina0MO9t
W1187afxWhCf5tm9cRTA3KSbNi0eqBICw574guVo1dEoBg5arJB0oqIgoCJO4+roOoZwEzudzvHi
wWHucJ4pVvTcu7fv0Ta9LEtbUKcDcxTiQ9w4NuWrLLmPa/JWwMmJbnCw9pqLw9BoEtYawVNOsWO1
WKvUAU0YdY+/hx389UOYBJ8DrzorFvfIvKP0cdtH7e3elA23ye++VEoJbH3CKtffRrUWyFl+4xfC
Ae7sQMwPdMASLawPUNQtckG6mf6tCteKn4JNIQuEVExnxIIK5XZ+QcO4Zne/OiwQAg4ei7Dai9eK
YXjmrW85xYb0S/Wd6vmXGNYc4yQXSSmwfzLK4OeaAN9kOUjjppRK7ZMlPHxJgUJCb1SnuWWY2+T8
ltjTnhbIanEiwu7gdYkgy++hEhLoT4xLt1TyobUOryyON/+izswYnmT+nrkxYoSvN5zCj6M0gC3h
tSuWlqQeff9eujinwNJuzShf4avl/KYsu7mXHnhhMnOjByDUp06hZlqImfkQlB34LHXguS3YZRHV
bPBrrX//s3+i2dnkB5HsSjwSYrE3tFRWt5zDU+01eYaz0ujt8F9mHrNUXWvIl389Ts+R+/Kb9M4Z
BUXHBQ8Ie9sdqBr9XJGXp2VgGxFyjsHs9IBVx+GQC36xQ1pf77Gj/RMyHseM5FosMB/9NRfmmiLN
tKCLKa+rKYLx7PEbq0aREuLaiGzJxx7vWhyIkXpqAaxD+Wpmhl/TbrluuCM2Woi6l6QE7ZWp99m6
Yap2h1F0QUKJM3X2X2FEoyj57P6VL8QZc4TM8+hxH9H4glO0ZCH03jjWwfVjZ6NOYw26LQ81bTTR
5O4nWHE4B8HVGTsuSMmvFFJD3viYavAF0ysRiB7FroILILzXiOCDZFxWYjRzrCoVl34DTOCfFUxc
tiIrkOxZ4oIYM1E3xXoXdZMCrKTBNpK0E/FnTh640s46lRHByxkrfCOYynKbgbmDpBSZkdZJsKkc
hj7ybv7aAc8gFQVhXNU1W/ZXz+u3Evs0c0zrXO30ycOafH/XsInynTscIF6vEY+RcX1/L+fk/Os7
StsIdMSnp/mfK8D8RV/YFJyAovlmqd5KmolrOL01W0V9amlApBIAMw5BrWAHjK2ayRWKj4TpEtc2
j6jpibkN+slJKAGXJf2aH+wZcBimeYleacI3NRzouMewxGFTzeUmyELZ4dHLw2nqYSoshUqbnVoE
lZgTBsIN6yQ4ypFGSFHLn4wFkznGY090MbPAeY7wafJM+ngvDUsaGWXVrrgBgr0O5prfOpF6WdP8
Bgm8jrV+odfASkopMUK3UHpeHhqVLpsiMoy5C6ogLgiNmVqZ9kaPHNx+kEWDnISKmp3wG0e8Wg9n
fnMeqWJCQPFEhogzstw5V9RNpcWbZRaUHhfAyXdDnAOh/3Mtx1lrScdgGW4d1xirg9t5jeHjgW3r
0LWwsMLGzCGfOoFD4UHY6RI63LN6gWWvLXIa0LdTJpzVnc7OVJJvY4tvAPQVNbSgtOyWRmBYmrCY
hH3+sfYN9LSVTqil+nU8NVuIbD341HiFShUmpxqe8zzoLNZMhh/CTEN7xkWkUzw2z6E9SXLqGZCn
5K/jlT9H3xcvZZFAAZ2bbXtVPls1ZCvRHO+ViVMqccg1o//7m+98KFtE35aWo0VN2eombJp9YZs1
HOuyFbXh8clGLxS0o9FIyyv9QFumrMHGBWe6Xua3VQCJFua+WSe3ZGtklqpLcWnVgn7VVzbv1Y/p
Bz27gK1GK/aaL9ewQ7s5SDS9EZzvG4KyEtdquIF1oVyG/KrAnZwLKp4SmcGXHJqpo91+KSBLS8lv
opfD6nu0BgGyUU4aXmjY+rbhpYNVR2DIxfccgBaLX9GVvk7GxaK3y2PWz8Gr0mAbySMLiTMWP7J2
trjsiGfGxLZ9yKdOXQaRAQckAc/HmgMnfGtNEkaPAaP5p4g90WQHVgL9XbOapTYQWGygkocgii/h
EceJpBLyxgDmFiQkiKwfyh5i11p8UPXGw1eAqSBzj/ovjuFGOpk4U9S4qSXafEZj8c+3VEyOwEKl
zTT54/P7teyxDOuim3e+Y8S9t0Yw7fPAEZJTBufmHFW8mTj8pcZTXSCWas8va5SD5JVYWfIrK3AE
CmRV+jxebOI//9vKeDm4c3SiGg7IZ/PDGSux6bSuJdjiDI8I/e0vKNH94w2yF7J+Gvdww3fY/TRS
NVywEoUhOBwig2mn9pSg5I8pVthw4Nhhre3O5jqUkvMhIGOJrf0mmt9/hVoDkgngpLVZM9XilkmL
hW/G9cizn3NzRtn4M7E5GSlyFCwRJQAb0sBQxAABlw7lvdwR0vIwhMPnV7YyhirxGgtPg28S8PqZ
0ftNoXm6czHfYF5yKqC/+2eO8B2L7pdfc+kqtf1n6CaBXy1Px43+RMLA17iZUMWHvVWlw2smD9Nx
We98QVRFecrTLKHHQCef98kxAXngOGSUhNZFnceULRmW+1BO/mTdgsnAzusu6Ojs+35injNrFADa
+X9M3OAC7LsXBtzEc/Xbm0TFOdhXewDSqqXuS82QNNooSHGkvFIsBTSdgHiDd3U24/NeRAYVGW8A
J9RMvSGiZuZcpIwdoADsXuWS5yHypMqP/0WHv71pLbbw16X6nypLqctRRogLbVk1tT6wPr2aZyM7
2ZWBtjY75l1kxJWCEyb5o+jHGyDQSVUK2Sy7IbT6/Sxr5ldkggIcBBLo5oUE4mqls8vgPzhcMaV5
OsTdV39jGTjI4BdhWk1XnNfp4X3eYoDxwIUO8GUFlKbO0En+TBELX5Tr36jnb0NVigVx81lPV6cH
NOSESTL3AfrXRgihbzKVYKyxpEwQYpmhSLwYW7V3nBMZa2B7Ho6Wig6RJnjfuA29wVbYxtsRDGyL
8WmlqHOZHMczn5Agqq7Bd8VVjNUOYx+8TI4I8I1hijt3bu56ME7Md0CYIfSo1K5+iauG0gcbnkz3
XJ03mL3hPPGMROxQjIP0X7Tvf2AhxT/bc22XtQIt87gqpafGivh9dufSno9CFkjAGtHutFjXvu0n
f+24AvO7dsKQDHPmFV9C/hV05pw2IKh/AIwWtIYf51klvC5ajgcr0kTZLhQT3mvX3fquFjbTVHnM
M/+b7CRP23FfvRsXS8DOQ9/7OaEwEh9Ga0pExn85iOJhALRdDNzNndqWw/zPYHuGsBCX1kpEhBPz
h2oFMFh+fS/l51nd3uhrOYc5iXGvjTuR4452yDDjS3q6XgqNSKR6Nr0+VTXQ2hP+EJalaITke8Fh
eBnDEi/w09W1qghW7y8dXAb4aOmjlkYpV3nYPDRPBr+NpNJSk8uB8sD8bZP3uElgkqEQeKtz8AQs
nfsbm8eND59JKjRIV8spx6CrcLAU3Fntef7LYJLXctvQ3QkjIbjHbG69F3i1moy+XK+EDmTKmqBc
i2AEnKCyFSlmnyu9TpWqkNVHBiA/340S2sh4f81Mr3mO+Gscq8NUJM395iQ2Y/fEn/sNy2Yl5jpa
whK8uqzAbgDMK4B4+1874DajZRCFgY5zYpigyDsNNCzn1tfIWojXM53frlBEeJBl4YwH51otD5uZ
Z9Dr+NU10chGqUgBj/629R7dL0tMBH/6Y7Ry5uAUSMJ+FOl6+Q+c2zCq+pr8LHasafULGuD6ao3e
m5GQ9fsz/vesU8jgKGxJrwPdSJHUnqP7TR6etI2FPYogC2EY5ayWskmgoulaHtGN1/8LBAQg2C/7
Yg0sGNdACpOCEftbBXMJkNJAQ6QNSIpnx1u3y03gmO6oG4PlAsRS7MwAio2bskezCOmB/IqF1Vom
rC0zM0AHCAEEtw+LNksTROZh+UXyroNLOJQLLHYvulkc1Bk7P3lOwqkbrxOwKY0HNHpKXa+7TNUG
6qKgW78tBfwXAjTUl9DLkCoa5HLESZ2kzT8jS9DZ+Ffuq/PY2re1j7LlMc//CIevkg1EZ4AxIH+h
eF4kpwhjr7xQtVl0n6V0QFX8Crm5RDzuFNHMqihZp2RqzOS7rLdHpu1bArEhUBdNFkvY/RUvcMOy
1gG606eHi5qHYw/oDXs3qc7OpW/kRbYagVR8vFuYrz5S7Gdua9DbBUh1T4M2Fu3TbVD3wz9BelpB
4Gl5z3gYi8Wx8jw5kbYQv5OBndAuPdLWUlpaTy94MjAFehj0ijY0MpGTXT8ix0kR/oK/pDo/V1lC
ZlKOcQ7WB4c4k+gg5+eI9lSR422UKIA6FGWFLSupnXKM4Uu3cFJoAI1MplnExw4fN1FDMlluhzo6
BVypM7LJkXLT2TOwEjq0WrvIVp3G+dJlPhrukUj6j4b2Ui8L5HpPMpjwWFuss5UZWQr7QkHAdhvZ
A/9pz6mLRvSYh9dJmnMv65DYvK4np4yz6ckpkoYQOahviDoSkQvi3mMEk6yr+svVVTRkDDWFtPLP
8nrSasm0hiV9KxLS1SOxBfvum8WYGFL0pNK7G8jJXYWZ0aP7vlHrJex8gIqkf3bqqVxjdmMGCpf+
lofcOdbHBAtvpMvUK3mAywDno41GNwLBY+8nqDbIykhomGMg1cHoZiqAsZMFt4dQedKKTAo5s/S9
RP7Y5AY6VNlLSqvaP81Gz+mfx2kY3Jc2UPrOI1WOW5twsN1uRg9dlYKmA9gI1Wogp6JPejEzzF6M
34X+KohbXW8Qmnn3jZbl1Ojgd0SweYzzQ51wS/NSXMZpM1IREY68q8WNC+2zFRnpzw8nuTBWXS9B
9Fv9CEiW33EIq0WOVyHvaiuKz32Vg43XzCVFuqgUcl1PhgRGv2C+92jPUTAkBPwGxxSx2rcfH3aZ
1qXPgmuvTQbDe4A6WayhKx34tulKDF+ciDRN+jWwtTcwOR5wqQ4/yGQb8v4LBjrKhio004fAlKcJ
AQKs6Ma+NFQPs9VJs72bWqO7fqwKHlKYOy4PsEKATgOyagcbbyKnNWHkk0lgsUSfNYyr8xQS5sJ3
ehSkfPQsbSpqX3KRZ+DGd3K3F9Mps2wRWs9KeUXZ0dMLg3VuxGdNzS5aLKKm1zXcOahgRS5imLee
sc+qy6JBmddQzL3KACCVhtnj3RdoZIpuSYhTxsD8ke9jAxYZh/+xP/XP1T+8QLSj85C3NRigAyaC
aTTUFzlIMP/Pjwl0tr4gh18aKlwt4kltEStpUDn54z2fEVcrHDJOSQe34LfW2FIuZhJyqgpIyJG6
S3ReuL86qZn8Wd44FbzhtpbNRCdQsW0nRETiIV2co8s9D19NGuWdpfW2AnVkMoHSE2QeK0L3DrEP
20Wm3PXat1H0MIkf3N4i5hACAwuON7mcmFzg37ueEm90j+J+eKM1DxXyHdQ+9QHrwInlOZSdEfDa
BuLDz+3kgcxI4zPsXgPRFEL+Xs7htUjCvaTz+FoIAOsYbeMQ/CpNLVHCJf6WwPqgYEgWIJY9jlFM
ucy1i21Vm+o/Hc2zz6NqgY3+LeYWEAlMLCprvmkYGRkm9T5kePXT5gOA8MiEyq+XCw2268YsTfLi
jMK5L6Z9Nmt2Qwln+1894+d525OLzbtQoXEq5+FJGXWUAYajUPeY/ji1OoWUj+3KPD8Su9ZCmEPJ
Mfm68Rth6pb9WSakibOMa0aKxgyXL5uC2a2H2Bzh0SHhcd1Wjx5zwYmYAjfbUuXwziMtVa0sQHgW
w4Xoyake+NqlJDPcoucLnM1LwJDftWZN4yTsHaAUNkpAbH5G/Y0QisOyY17a2ffbK+iDFbmyM5fq
L3TT+gYDNVj9H/pPsYolZoqT6cSwsA7kcf+UWfjkqsTUkwdP1POkUOnDnZnwRa70O8pKlnmyEIpN
jC068/5ilA1gMPuF67yfUtxNHEkqcFcS2+IOvE2wLC10L6QWyO8eGUe3uM3rY0Pn9C80ogsYvu6f
5yOnDff27ArxS8TW/LRX87R3+JjTeThU1jgYIKtTwWmPfFm9EGFJAwyLfLYhysM+qMH68cgNKTys
fBt3przjUMLFx0pvJqrs4FkJM6Ids72eLRe0UcrlXP3SBlPmhkqxgDfgEGACm7He+ahET2EF5XHU
u+MfnTfMMBGbZ4dUzc6xiqTQzcCktQUsz7AjkV5Z7dbSxzVNDViDnAp2R2g0A6aG7DH0r4wqxJ5z
wDKyqIgQiP0h+H36b8F+HNxV2qeluJwW1eh1UA5G3tZyrysC8vnLwQMGkmv7UfYQ0ehBtmyw7Kpe
npvk2PF7tCq4b9hSl4OtZGJxQQxuboss5zlgb8C9OiFzb+UP8ozzyPDLaCzrr5LaCT06sa1NiLOQ
5oz0QdwC34H5FbXkmdDHTEGAFjPnK354sTWJyQF/IWGFg/vuxA40VEHo5ckL8S75+MC/c3y+5Pwu
S1JrUplDQXEOwOLhNb+lweDb8y9cE4W9cP7Z6IdeJzgNKB5dgRcNMT0PWjQYoHUwilJKLmFynJHY
Agwx/4MD2O799kCKg+t/4cGnPPtEkpPz5PHp800kk8yUdjZAdzHhApCz17DfDf/geCZONsZM67u3
eVh8Q+lQHZVgbJTTPTe98WpthSVrRm5KDBa3CIwvECRxctFx/qVOoNlWa0cx2dEi8eIVVyhj0X/D
526du2NpkPq+s/fd21SDQxsaXanHM/IcoPaPsgUdpTAGfzuVdBC40HKQC9bIOx0YgtCqMHn2nfa/
WWg34sS/GmHuOLLRTZKF/iSC4b9GCcDIbZQjP5JU1TbSKuV1xzhJZLl91mGM1uNW0pwaWq988BeH
62TD07Bzc1KDcvtN0oDWw8LVV5T53tpBDfp2b5W0pIEzjNpIqcHMOAp6l/5V+FOtSH+PRitqzI06
uTvhINXIacY38S0sYhZi7Fk0QxCB2i7tshbX0guHPLJzhDjX4bJOjmSHQRs94qFQAdbJBySqQU9L
3lXLmdS9V04IcZBhvBUu53dwCGuxp0geubL+hHYBVbOIZ+wSuO0fU8R04GVSX6C3u+J9nZrQO4vc
afwy/GnBeFOPoQ6o23PexrGabkhURNP0bRUDCshAIfqtGPfC6eCEBooBHp3oV4JiaXzplndxLkNE
rqBZkyL0mX/f1qUHGwmi8CpVUM+QHi6syy6Dy4A/IlUIp52LHO7pJOmKglR+lrx5a8A874xUZbZd
l+dNIkCt422QNTS1s1Lyj3Yo5G8VeJg0JUSZHSvtZFh/R7rDKS9eNvtHYIyRgt9J5RK973W9iEUa
pFvT27YuSPU6gXuKQ3nN+WZmwgklCV32+xstr7m/aRZ5VJdIckzKXtSo3jgbmVoglQrniKuYQETt
bNkpv1LfJfzd2T6fdtBezQqRZvGcpboCDEhl/L8h0LzxuQGjC+SG2F1yysJy84dGTcZlXvNyLPq+
2cq95vCZgoQCjAejGO7aANBDW/dkQWmivfeh00d+cfLVYpccOIXijVxzeAHqp0szztxKZPDIWarq
dnHqjQXKDhfpKorHAucRi9p3rJoLW5O0wyB9x8TWJf8HaMUOHENlaSsBXsMp1mUdZt6hU86JXG4L
BFKi7+HIG763xzQZmV+qFYT6ZOSOiQydypUZEKrEd/j/3UnhlApS6+ciPMz6yOluNH8KKV+J9EYe
UNbIQDrX99CTZWKC0fcpVRpq2N5WmZKQN0SoN7triHt1lXTvihAOjGYPednHF8bMnX0VcPaCmfmu
A/IigffHwQTmEzoteOGtumpT7l6Jx904tH//qk8QXlmTEcJW5BVwP2h1sTWvdYIIAurOPQDHhBru
be7VSMcOZDC/jjrkWtcvqDkEwXqTsrSPq8hJ6oqCGox34hAwN/oCcluuCBJ2yIDN3BuszvMc0ABB
T3CtuJ2G5c2tGQR7ZDVFokO9rp+1qJvSATH0axfyheSOMSP8zjLzM7r+yRoHpx39TFdW7mibeQ6K
tuNkF47y+gdsxaPCmyPAuhe/ZevRiKFrD5cz2ks+p3hauOiHPxYHTGdPulAxvpV5iErUlBXwxSiY
Lgsw2oMQNMtdaevwbMZ1DarQ71vnuVuoXv4IZ4mTc+adS+JDTpOxafT6STcim9eWn9H+2VJM5o13
qIqD7/eQuPMwrAnclVXiJ32SdTbANRK/6NqylBeLaTIo0EcU8VDuMZ4nCB8+It7zPOBim6QkUk6j
q0GVElprdUnFGehHuU3FfulQJN/wIhZ51BnS4hBww2ChUvr9+LPozUrmi5MiKTLa8M5pluIvgFdu
pOUAiYQRhVdaXYku3Pgll0Y21ALWXdT3rUeUB5GemAAhahJe0vkMue8w8vL6q46VXCdz2aP6ukWz
RyH/uV5bQtKebErEpjNbGMu2Q8Cep6JVcill1k8trtItg5HgMy1ZMPnu+oO7NqAioAByX/xuGnwO
mckBTzZ8x00I3elnD8knOauqsvM2y48Xdp0uMrcNshuZJg0Exz6sb3iw5gXQdeoCBizUKZzJYSlX
a8JeQnCr+lh4t/Aqo3wCVxvHiyqpvDDkhf3ZVcrXX/C10Owv7eEvxxoNk4GvoIUVbcd+NI02D19S
+hHErT4BPIdAa0Uv+S63yo12FUxwHLFPLNaCnjrZcilqyzz6zFRuye6c1/OxSafymwpiON9H6lGn
KHdnDjk5doEOlhpv+QMx0T3n2hUynaHLCOkmjzoRIJSSMCd9otykCXed7ZwG4bVtZF9rGeHvdv6f
ur0p0rv0qzuEscqgOkRDLagOJObn5CCesKZnV/b3Vx9n9UBjj66lDWH2KBydohkgBztldHHqRRVQ
TzQywWj6+iXEKzHENY9cNP5Kpmbigr80krxWCE8jVAZiL1OzHNzapg72tS53AVj3GMpyPHgv+geQ
7dS0RMOlh2lfQw+ttNEGUlxmBfJ9Ok41KgIXNA0ze9gdpf47HueRtd6RxnrYaRdT7EMvIQQsVWzW
WqCHR7XZR++kl47HTHa6bAhwHwV8RayArbDPFE0zydqi9U69Z1yGEH8vM6fCRqQONVuLQXWmhZVp
IfmM88f5zEjNEhPQNmQW78VKaN0dQpHdWieE9nghPlPkJIAy0FbR6O9BwGkCj2MItAzCQM0UW7oA
np1IaB/OntgY4710+KoEOtp77+GDNfltpRy3OII8BgQ/DLdeAcsMM1pfcnr1FFAX7JuTewNG4h24
ro7YqVeQi9rSJW5wr58u8GCKF81DrzfwjaBgi3VsBZw4L9gFLxusJhNW7CRnRsrJYfqJ29rPhec2
T/qcrwoR/0SpWe9yWlxOPf6pzhxo0uEqcOm3o081PQn2AOSS5Q3jsfjGwLsFlQ+f1e3u5xnLpcMM
lZIfrrlKy1pXkQtu7JYg7pNmy6KW10Lb2+fG7inUz5XW5wAxAwcz3kfafDAq6OYdxuXoDmCKKJi0
PNomWnyaTulcxA3357d2YehRTgPogSsNj07yteQFnr8YcCr2nC6thoPRUnaFfid9VwyxHbbYccBz
uIqkIJ2Q0en0feUZPDiVRGpZToqOI2WiLqU0D4cO1DUyyaD3xZakeTwyL7SsazfQfY7EARWyf5lc
aAmKdSbxa2oHMlr2fHQRkv4/OsON6BFOpREM/+q/bozlLSMo7Euzj4AxTSC302ZJNjaxwqHwRcIr
k/FDaUrFTJ+CCpF7iJs5G2CnihrJR3I4vJlB2fo8wwDQMoOTDX7MLwuIH2CuvM5+XnyaPxRvfnxz
8HFJs9baulilIG0OTjq6SPwlHG3UGQ/FFdv8QgLP2ep5YwOsnA9IoECrZPdtKmA5dNspz6261RRw
ItaswXK9gQ5mbThxp8mFA+p+V8BjxrEvhIJVnj1qbnlcUiJyfph5gqPnDQQZvhOs40Txccah9vo7
Si2apDCv0InPR6rr4ni2fSEfhY7UNEdl2za4qv8EoY3EMrVkFI+jEvywcTLrgqAlZJ7FQMGfD0NY
ghzGXVkrReaar+a/bagMhq8b4ecMS451Ytx+OTQ4b612sTbSVi6ppBWuXVE7oO2YPhZ1i9ClfgIs
l5cTjRCQpGoi2hPSNX5AH6zlAzycmrDzvOl6tUnVZfbiWn/JbpudvpXxMJ2ll7IY9fx0XnejSBXY
V+h4ez2nKYoSf4r3pcflpWF1rQ48H/BWpieYHSbbqt98G5fSwN6JuFK6nJhByVycT7u5VHtz4WJs
T94OcDDfKbAbtuOSPplQiSXKnVK2w/CwDJcuFRcWGRf1hG/uUQubCAZLJNHRIRnXVAsxu9Ao5hYZ
O0LXA9Y/bCldBP7R8RwJiUXwLMDE68OP3qq/t0U/83SkEtjr0zq1YaIQnyxtmoKk3cyZhtoR3EWZ
k1kXX8et0hW/SSCPQsLdrSGApAF7JORUH5NjB0NQDX1dsLXmZ32whIaQpTQTKGot05MVVdyaFdiG
yNhWg1kv6Gszvg5L3Qpkiekj7znBreZkUhZXR5/rddK8ojH3HA2cET1CGrUTyFIPTmuCOguMiEho
6HaJAJF5AVPw3/Xpq+1gQ30BlrkEAV4Q2JP6wk+V2p1ft3VGnRY4By3GW1XlLfi7cyyHcxBaPiW5
lfMky0BEPSqTjDz8UcmHE4GF/h0NgX4J9H7f+lRgrHbXrkdNRbnLQN8EY35UGwLcfttDQpJt2sBd
FD6pLqbxKl+eCauXwRzuE7tAjvJKiKfslznOzQh5HZd/QIHpe1ExVzhcsqKa7PCuE6sqnvSJvobo
hv9j4tZ3Dn5ot5n98PX8Qs/OtCKzcyLK2qT5qerfJDOutGE9DJlaBqB0DFI1ykByeyA6Kk8eVCBR
xqATvIcGO3sHYyD4eYP4u+yuGkV3aXmPFpoy0FoX6AINFF1Wio3nkmaMnQpmZtt4q4kGjwXBj1BZ
DjkpHh0LueHmzX+4DkxSwBswvzIFDK34XvijHtcOVuiKoXdacpmCpAvRxmMu6PrubAEkaievXYyc
X4H1tjkfNKs9jWuumGzYmcZs7PMLjZZJo1KZk6gNTK5JfUyb3BOWJZ62iywMsC/TFTQAJCg4ElkT
nfXQzVYUiKPMMespyT7v5cop4/oOGwkP/kQoSwUyP4fS6tPEuZVRVSQqbOIHWMa//j4IrsOVU6Qe
fDPmPQenEApvBgSrF8CvBg46q93jEZGzZllutprSOxnXoK8yK27xiw7NMNa51yDAe3OE3qYhhm6C
xUNK4J1tYz4Zx46dAlZK3yFMpDUbv4h+uDQteGHbXSPJreQE2S5/tDsoN2mAR2rkfdk2wgu2XG4H
v3+Vw5aTqFdvwG7beRJXjSzQWKXnonD+kf9srT+SYDFiqEm/fsVygoPc8XElUS9W1BewR4R5EpFm
7XUpAdOxMJFG8BPQ/uEwpM3lszbSjS421LT7F0irdQUphpy9KMKe3QJj0jdfIP6c5UWjI9OkEnri
vo7/ULTx81P8ZqfmQNGDr1OydlY/ZL0L+xRp+6Up/+HNzNOzv73PDd9G1B/gHF2RR2LI6c991L0U
8fC0/tg19pboUQNi1H+c2dkF78CnVmIVjz3U/D30pDDufsiysLsSZAxU0yNtFIVIileIF36qnBYg
h76oVr9d3nqbQsp35TZW/o93CDBLKx1s/RyX1rBuLFnjMGF6Bw9c279FErUJrU8gTtBNxe02UUEw
e2o3w1NvJAlLMpnfoJKxe68n9Y52h7V8BgMSpsWuC8HNpwCizne3AaPlmAy4jUPWZVu2bogToZyH
sA3H6Nx2dVCUYXFBy9hFLz+OXKN+Bj/2xRrk5RaFZNr6j0V4Ba8X2ve2kKbj15W74497tk+NM1zQ
N7zQh/C6PtbYyqRbDMi1wdJMyVBohh3sc5PWWDzGdqWimqv1YjK9zBM5r0azXU4ZmRKHFRUAOhdh
QQDbsjBjKUDxD/8Wv+SreUfZSjb83nxKizQ5iff4VnWGs8XFraE3NTRO1kPj3TBalh5tjJypwJza
vZK3+OECmVsbvm3VHg763/IBbKie9TjR02kmQCrnoQjzwyVc4GMnJe9x539664qDq0owi+j+0xnR
oO/8VpSOJBCN3M8YDr896/lz3lCYEOGeB4xgHyU4koWV6gfUXGjHIDQ+qoOHFjrAE5ndp7/B66ve
S8HH1SKGEpjYFsGdezV+x2hYjIWR71nQ0x+sfrLoTv/UmTMarRf6Z4itXP7ezNreUWxgSQlS7g/p
WpGowXCAYXE2WUGRdH8YpPBsbl0HItshmu9eHhoyZe4cf2IsrU5YA/XJ4dXbGjXwU2cf2EdXeIaO
y2DHdDP8gpMSOkcfrGC0Zatw8vMZ/WeRGRCK1U6T8LZ+pZrhdTRdhXeqkcMQDwoEi0jpjSiJsWqE
ZRIr2TxgKqmwvVq15kReRtOREa00Nszr5ATh2X7EewkJpTSLALOP4Hr+sOSnDqoJvHYfqnk+v6hB
A59AUVsEyDSaAg3LPu1jzLl/X9okQJkqfdZGBadL4oX6uJuw6HHamCgOu24ihOIs55rJmRcucBvJ
5BnhLmTq2MoRaidqV1yR6K/KR6781ZLL1Na2KZuXYyefVBJ73PeEhtWPg+PB4d0xLbPbum0TE24Y
pd5KgcpaogcsG47bR05wvSwiaTQwetIsdCm/ubaxb2J+aqZlPQxLNjMCQ1hKtpDRqxJOXinVbnB7
go0HGMT1/3zsj74dYUAkZuKgSumk4Pdw41Ot8u9rBF7+qKnHoSpNpK+uHqDg2nqwJIkYFaJkG5C0
ps33cWVEr8tfEFNvq6MEiTdAgDR5UeVGcUrlnaDU43dzHA7QoJLqCcC9OKkKHr5k2NEXeCywVpA1
a+ZaIusXQR/Ju3ADO1FfzgNujFBZCdRuj3RSveE8haEmohaymgGG1I+g/dvTTRjRbFjERbpJSntD
UXUAYSpg4wu+wQPvGuJ13EreWxlFhlYW8OX7xfH7Ai13TG969g7dUnFsOSLPyDzgGSA9iTf2PT7w
/Q4G8VDjTg+Zxwo6tSOELn1uwTBriOparZsix/jgAAgTQYsIUP0oF96RAEUDcmUjB5UjJ8jSiy7b
727pGRgdxExOdexR77+WxS/2UFS76/quMaSJsJn1yzZGfLi1kPs/1V6NBNRzwrwLgtYQjqdUb3r8
145qaDFtHSiRiMoarS7+kV/B8amFOmjUXV8OOamPibZsi6/mtTaVmusiC+wylrHV3FTj1K2jC6iP
NrG6bM7MUd43+/JLnHIeB42TGO9ZU+gLe1pN4LRHfz/rKngboZNnCWpNJT22vAv/VNuf1qyDQUaP
HNwem6VpPMo0kAFeAvoFDcrY3x3iR38c7Be0lqKih/juVBGUWswYNJGv2FavAIU6ckSiXmSTghWS
dVV/l5ZRAXF/OLjFzLnd/zW+AiQLX1PTN+vWYAkELbvw5NfnZfEzMFXjzkGXihBLb5mAvXllkAbb
Rpn8n6zPMRc8W3YIY7Hv2Z+Oo9m5NhdWP3eIZhkDE2zOrClfsfXTgw/kYlNUvilPsZ8gNBC/CWSI
irM/KRLbvzX7g42Padet8TgaA5tTg+6+8K17xKh+dVXpDISwX2y2bF8obXOF2I0kiFz7PFABuf3O
vrIyYk+jH7QeaVO2aKfuJerauNi/zAyDxQ8MP6vt/iUYcXwlriSSGSyOOucZskRzwY3HnSG/nGSO
O1UbOKSgWr59OYnekfTNjLhkDm0iayGB6GcPTxpNlNIyOhrF6Sekh4gu2MYQolSis0t1WMe8qBw4
MjdejegHtiDiPOIu2oLc6U6NICsypOp2cLLaJdfECA4PbqxgDnmY4GAdGXNIFTcbfbPKnRq2L6Z6
BLnXuotzhSYJoynfHW/GCin+mhWzzFVe3gqXnESsnYPXj3F3NV11dy3Cl79pUs00Efjdj3LMbx9h
Ab+1AeXIir4a3LWkrXmwQwQOnS9FxjONj6PD1LStfdR1c9HS0WGQ7Au7k2JcsxZs8BuTu+DMeKSf
KzvMVV6rsGrEvdyw3ouDArsf41zVl5uWVu8uNzB3oaG8ya2q8dT6NnLxTUgcJ798YkMRKXEDNqQJ
0QxOau5WiRjnwYe6S+3Z7AJcnp0+FEz/D2LlLAEZB/Wlt58I7I33KpCYENEP8rB9yeWJUZYIHkpT
WTOe1mnyKouA1OlwbwRmRgAVKkYEVH+qgYm5IDtKClitcbUMUYGD90vf9eStqDI45xy8Jh1z1f1D
6uEPuVgszaihyVgu1z3bJZazVFSXH/nmWt1qI5Ud6p6lo/ecPyhen0kFB9tex7rWGwruJQm+HCkW
9P8yDtEg6KH5c/1497uGEAeYn9qpGL86gTFsUffSOhCIs3RD+P3nddDJbHRmD9goxjJeNjlCTzN7
SPTGnlPyPr0ysMvtjFKjoOTDVY6B0ROnIIj32d5bN9KZroOA37NcM4ohHVtH0Dzl1jjUJGotjD/+
K+oDHv7sxiEfNe/cQpYot/G5oIrOWZPL36Hfuro8VI8Mm2qF/K8g58F3fzXj6rQixNUqCKDjF/cM
s1U2titM62gm1eVfVcljdPIbMpGd/Mg3/g5Rblfj27t4pdEjUUMVhqF7ZeQfsymx2bRL64wV7ptD
gF86CQXQ05Q8qiXvXhWL2SU8kDuxrUYzCCcB1rwWJIVI9IFUrNR/Ta9iAzqu7LCskkuthA3tJOjJ
LjjmfGcSEArux2fNbkld8OIrbfcjpJXTSaaMBNThGGI08kqKtyeFZuxRssOtcnE/l7Od2rXQmv7L
tmryZ42kK8e1TWMOPLZhkSn2IypaeMuFKqg7Ft+4XTNdcMWI5wIu0Tvl2oxjCMT+dAzM6rFsXt5K
/QtG5TYV+u1CC+I0sRDTLIi3k35VYV8lRoV0sVqdzQ9TTuhhHs6+9GEeBFR71GtWlHqtCYLcb5f+
Cjon/oHT2T8dpHyLBmVGEcvex3WU17KdDlfzHEE2sN4MVwWEmzD9vrsEuhf/mY3hQth4ol1MGBj1
SnYbUWPl4ev5hyv4kL+vkAtMEUJnXbNrClOerzhk/wGO2eG31aUNVBVM6ZMehHVNDBNqbzUnNBQF
VurPmZTD7PZRxuFSxOBdKi53m/whTBINkGrwMHG0Pq4g3UnrXHqZE0g9zwmjtrqn98vnIb4bznuI
9S8pHbIX8cslQWoSJ8XUqgY6POHIeKUJJSOzoIJ6efxAyi4RWKLcfbvqDzzjQwO2B5tCB/N6UF/W
4QR/+O/8toj2IfA40hLiiPGs2lVCTx25DjPwb+K2FP/ehGYMl9f6tBbwhTnBJuCouEmnkKkvn3Yo
bo/m0EIv4AY6f5BgXkVuHKgY2i7xnoyGsd9u5Xi0kJH/tJkEHBgG1OqpBUQ6RNHZnz7Ei0ZGmDaW
dn/zK9X3APfjSiy0hG6doPmxf5LZ65exDquSnbNcpNJUVGPoaPph2yeR2PaXoYWLU5Pi3njuGNSA
pYw4jmHR3c7GIiDUuaynJ+dd/vzZ4GEPT1O78T70NyLinRNLLHiGWmB3Zx3PADMx7crxfK1Gwdjh
rb8Rfz8uTHa3AoK96qFDN+WypfeKGeiA38rnLG1mYLRnbthl0Jlqo/9PkXzSDwqnQ0drAj7bmNoT
mKPpWbpU2FHDnPDVj57TR1IZt3J6nVjf9H+L9fip4IA8Wob1zsnud+aqXRmuVrpYb5f0hT+AwRhW
4hZDrd95a36bxkNTYubZWT7jkz92RQUuUoR+9q0Rb9qWOPQvhu6KRNEXFkcMimdwPctXuzDZVYm+
CxXxUZlT4i0zaDGhCeVOYgq4idtNDlHeirS52oYf87wBTnLm1YZA0lc5zBwf8HvOC27JNdzLXgBH
GCF1kf5LWIOEMR05CwoMaqxxQFYg7ZxAXsdXfrYKw63/RX8ygfOX2z0gAuDXDF/YipKZgnERR5Sl
O16TDQFtub0e8PvdFOLeqMUy5gIKLgitTH1C2hJ1t5mNuTAE3BFzwdE2wvVBnI2PN+UjP0i0wBHB
k7P1FYAa3OcZxvJYQQ/lWzx4L5i2jRRpRV10TA5jZQNdwiGUvom0jzTjQm4bAUEJo2kyvn4k1w7g
VM3aVjIy9tRjkbV01crJFQZu2LSCfHundwrZipG9TANWqIDqTmgwjJR43JEuTHcmFjIFgBphfzGe
Rpz+8Qun5xPnvaczq1czq/brWmwXYhletNYMy6K8HAKs+ldOJ15pG0PrjTika6HRhQj4PWiEYmYU
RjAtuJdaeybMz8Q83LiabxBCT11dqbfEMJoqQk22/3nuv6VMRZHOBXICByhCQgmAyOITeP3dLWfl
PQt0W2lYtej06W5PE3M3iGM69OK8AUQQurSsnx8gFgU1IkLbC5jBdupWPghcdXCVP6TVomgGBd5H
MhJ4h63ELmVlUOFf66scvL/ey3A+zz5PcTHH4He8biWqZsYek9t1lpz9vVG6iMlVA50VQ93pHgjA
St8ISduzrjxPDqnNBVlorepELS9QaINrS+jMV+Hu59Hosm3lCjZ/FoDdlo7+hxAf1DtEqARKOqKR
H2jNt64ChuSGYvT9rIOnJH1yGlkVHTSRjVZ2a9S8YSt9M+3yXysZxcNKN4uY1rotU5dXc/Kr/tcn
FOtvQc0LnLQt/Rxufh+zFqrxha9IOTN2nahIjYkf7aoCbCpnxf8sCWwxv3CIPlclBkR0B5UygwEg
NZKCu576lK+HMBeRAy/EKaqkWw80Jf2W7GK+vNJYHaCJQVCiI+9+k4FZvTeXvlp2KdigVRRdXKtP
hE/fIGWcf8VEhwKQ0Z16fBZeMOapZnW6Yce62SQZpruk/wzBrI/s+8szDVGdhu3UwPXg278N0s7j
0ohI+0jEZ2S5LiaJuyczxPmSgseE4BvrwBnZfFAdrh/+Lgj2XXbgO0AmqeTpAQxVV6GC3TOEWAYe
R1i4X73n3LA/0eV6eRSgHHL7NoHjs2/G3rq8PWAzQt9tekWK8QSRaKghwwkLyi/EHYXK/lmQRfTU
z+Dr+UzCYAMmzdsUdR8traMd/NixEsHw4QfxF/W60k6UWnrA9bSsWOqw98U90FOMyc8aVxv3o5lg
ORQjh1y+5OzsTvWQHbEM0dsG/HALKmEcV/YfZkhAnJ01SJH/mIQUvTTZoWsTbCg1rHnmESzc7xMc
fziraKHIONmq9hfTjGrkVG0LLwFtCJwrQ6n5T4pw7pS5CMEN8kJZl/k8mbapbqyIiBgIVQJBg8GQ
nPdbhlvOukYftJX6FMnCSH/RqT0dnrweVz0FywW7Us0ALUNBBT019WlmCxYIQXovu0quGJX41DVm
icxqBYpa/ZIm9tn4l3HN31ZHRU5kHHPWYMxYtoHtgHJ7M62kTbbzgEge3da34+xHitT8/vY5QK+5
54HSknisIqrVodEhB3bvhpe0XwqWUbZdNiJv3sUBOWufnMJfuJBgpfiUZNzbjnHiyQ+OJggajTnk
0pZb3NAwegOGRoeP2hlj9TJ5r205tj0J5CYomoS0+/NccNkzs7/SjENv+BxZGyjLBzIqxUud+5u7
qNjJ+8g09TB4ZQx/ocb90nDguqhw4Ix+O+P1K2rH/HQgMfKqtkRhKhgLEtjcTrZHoCLPd8JtZd8n
AB6dUWAh309txWPEUmsNHeKyq9aZ8fkKtLWNbHumU5/lmox/CfzeBofxMf8GsndtrUHyj4ed92W/
7e1khmx5ujL1Ni1lP9XsiAbhtzuw8ZNWaQ2Bw6X4TO/GiS8fZImmXFqlqhK2CFSuQBhjQJfQWI4W
FOs9MRyVFrb5TVTgiw8w/SVWbMBFbXJ0FbWEQqdgbu2oMuOFz8/gy+jzwH8LFvCCvsFtz3ACOefK
ecgFdxLZ82jseWWAOxfXB2mZwrG5ubftFbnT8Gh7WuGvLYL/wC2SEv7gHv7VeXrYYoFSiTo1TOi0
KoIutkdBK5aBsBo057nowgEgESbFbf/wznDHjwRGOSAlBCAMHRzSqFE7wu6N/DNRwRNDZXCwhs3O
qotnUZrOP1Koi9C1Q3kmXp16klA8wUE3iwrGSHKHsq5acYFVUGsVrTI6bo9+uGfXXIkyxnHJIdFN
j2zMUyVuHnzyTctqvsqR3fiMZiRDkvr6i+EJs0WYKfkW6NNxwjM2JD6yqoUDQBu9WDBD8yUCy6Fk
KMDGaG9YELW1op7bRj8egNPSKBwNyOkbPaI0uqLTR0+DiLxBLglXugeRzBn8/vfN2vfH4ZQXgaOT
++QhvCeaLF3NwWN1kuorb32Du3qIyeNkpyw1F9IIP2vFzOSk1AH6Up7hRtqKlmFVeHTYjgzclyqA
h6wsvT7RnQB2VHRvfpDAZJhBU6kEuOB/vM7IzjadpM4hAAUjIJPyYzYmTIQ3jKUeHnE561Ssc5IX
OTRH4VGUI7vDVe1wQkNFzr54i44oCULNWW1a3Ty/nO+mqk4l9n3WxAAAw1oZcu0AQOD1jsXHtZ64
1lY8Jinhm2UURYLeJ0omHzlqGU8zr0pP19pyM/WqygpTNJCTxI4ByAon7uiBAlXbMmUHV6lDDBPN
VL4YzLwD2oEyBvGBI7YjZ0FpU8PqFVXBR012pf1bW5l+Z0Cug5i/+VcUWQVeXDcVCCBlNNFf1Zw3
A79DIhAVoavn1dLgKwjgiYQq+2+Mw0keyectLonuRT8O5/M77J91/P2xzKcu7ywba8NX1/ttB9ac
VUQ8oJwJUY0wf50EEY5PimjFc5WaaEUo/0B5fIuiwewrSUF7G7u1X75e0LHgAVvhjgl5TF0nIhWB
7pyqBh4iIJa4eKkrPJ89C6SAvNDfZIzuheCKEQiz7HI7/emktLIOpzPISxHKwohGQuaLldqXrh32
RyhHa2ztz0PU29mimFhR5TS2zR6RvdbndFNjlqMnMnsHRIiby98KhrhoSXsm7c8eVbf1F9PJ78m6
1JervSC9D/pzi2/EG3lhh3iY2ZoRbAMywqi1Ay5SkzrOV0+HOsqOhQVQgpa7ZdLlojiGmNewRAND
UlcK+iFlPHCw65Ne+WND7JakLLj2PzGWhkl80LM4ON5VlwKZRCkd6lVCQ+c9VEMjmJUIuD/aP35T
TMfa7PlEdsQmieYy6QaOrTadyw0L6qovyBkEjJL9RBILXQ4C6oGgqOpV4cB9T0Bc4rCmB2ELN5RJ
eUEcagL84Z3citYFH09DMsTRvfkbxgQWVmug07kYHG4H4LZ0A9SEWiVItS+pELLbtetjmJ+7ez/P
HK0nCFD5QViwQbofno+n3Ph9YdvtV+U8OWP0iS9qxEEjj2ZCpCj/XpakpuMV3WS5D6rPuvE9Frw6
fZlOEF6aNDUlyAzpKXBYilm77O2pdWJ62Z0ifKlsqmsblUPKbfgRCdiPORSRyIbyGorb0pTcq8vX
l7KAOS+unzQuGDhXhM7aAd0jLIXDW+fLUwNF7UDIqXENFrCH1+ICloLgiUozFc4oSUTaanckkJ3O
yUmlN/muJ0U3RqSmY8S5DwG8LAVlWlJJQ/ty81EuBWhyoVJVWICNPRQatxLx89j55OT/T4cXX2gt
WhGnvBLAQGMsZIuQ0HVdRqB/P2ati2/x2fWMNOJc7LfiQ5dxaCzqySerP9ueltafhEEZUijNLMi1
lG+d0yR5Njp1wAkpeOhQVjiAkgk/y/bVp8EChUpi6ot+8wiANbNjjS3uy2vLSx7qxXQ+mg4RT/Dg
3EdkN96mOGQSomQMbkqZPSAcmIoPc1XTRVH6EEWCvmGTkkY/ct86h5iZ3Z6CDiKc8pXVysZdEDFA
uzvs5D8JmyJqYofe8z+6PygpuKc3ma4AewW2YjkOIyDLhBzuh5Lwr5N8Z4eRE0RVUaDQVqJ+1ebm
0oEpwqlOU0Kp3CT9Vu7ne+bbMIteycLE9gXt5iDTAy2RPe1S61Jr260kypzYFiAIk+p83XqkBSS7
rOQkY9nqWWWHBLIQGSozaefnGUn13N4vVdx9nKjwuElPL0KNXyMD9UMU9MrCWpP1U9k/JOH6QwFE
qb2s2LGIZHUlNAbvsIrn1dS/dNv1AGMEkg2Wu/JG2GHL2K44028SZEtwaDDeb7Ka7Fj1zW8vsXq0
Ka8gUv2xbK9xjrK+nsYbJWxOBCdYah5JTpjHH29keCbRzxobv5V2hjJ2lG2EYkuiIhvUX7LOP0kv
VrAwlcRiDnCxMrxvw4Jt7/SxcdMYg6TczSn13wDxmny2w103nrlEunTQtJE/IjGpWwNX4B9asMxU
WfVtIM4BUMhjTBtd+rlnjYZagpuCWsT4oj+gty5a5S65uO/x/K1ME1CVmnz0GgDIr2OBPBgW79Wx
k/iGfXsU4IFuPQCX3CJ2T0PahFu0fQC55B3dETzfwWw9wFXBmNaEm4XvciZjJ9aFv9oLMAPP+zzK
oz2qFNCFWTyZVBBKzzZWIK/eVdu60pTbu20hwKSJv/TCvHFnOyaHj2aDBnL+i71oP4j2eRwilHq8
Avkx8Dl9aFjoRn6XsXbJRkBmCwTNd6ZAsRr1Is2ZQ8sEFF2wZTWMGsU2GqAIVXTY3y/yuEiWQwvp
zQn9Y/8f2L996/7E2uJUUUF/4bKYUuYW/adee3X5fvWZ6PiwKoCEGnM1+fHsqVNXmtYIftrWrbDx
tLkfP1boJtysvX26H1v8HGsQffHQZZvV7PSxJmEl4nesAlm0x9WuzZA7KhEQQk8uwDSWr+0eFM5x
w/5ytMwgGnuRqnpH/7rh1WWbgnhWgsDM4JUSf9q2VzxPGJ9uMWtBkTWsXeE0UhT2MDz4L2bRt3H0
J5FvOP68PgXXcjU3Wv4RJINgNv/DaHNdl6PaAsOqhMEjS8hQKu8OnQu5nJlz/RKEj/kdiRAIeLCk
lUBCwWfk9z5mSsm7kHsfVhfDq/Mom0c/V5+5UGcXAFXbGCRuvlA0qqitK5hbLVqR+ogUDqjlM6QF
6HLHhucpj8Fq6eAU6cTX6ryj1jHU9AJ5pIoQ2ZjhzBGfTKXTia7AAOVJFtQIHaf8rRDUh7Z+s38H
b47FiXahOO9sBxER1vME8B3c825nDxGDRmH0Ul5uqLHzFZ8FnFf6flYy+UGuPQoU0lSJ8mriWv19
day743VJZPCXSc05ixrkCYx+GNEHR4tNNdoa35j3EI7IgWXkUicD5YscSOXKEuXBjEfqqfWjy5/c
JoTCOysTu1JjHmXWfMg7td3ISQkvHCAE86mrxy8mV7v/jkt4LdUiLf5PwSrPF/MUcX+3mi9A65Dl
atin8fLPuYWXXdEzDUH/M3+kd977Mu2WvCzAkLOrDEoL7vxYaeKqPnKhoZTXbItZaAxLU2g6AlWi
iclWcrvpCHP7WCojtz/RbqOtdqlehZ33N6DAF2t6sWl8mfT3ebU6FoYy/HE9pcqXHwPsy5zYU9Ry
+f+GyqKvGXMqjLMmGevsyF7otslwO2YkGWWbgIIuClZJH8m+uFsLBzyJlAhc+esHHk/37Z6KfbkV
qnIgz/KTBw3rhqkT8PWjH4vQ/ZyPKNNsP9iDRrsicidrNY8OVWG2RlYYHgXgyVr++xRpy1QMNe2z
yh6zr0tTi0B5wKFoJptKSQAMr9onYXvkt2VAiar7mTyYHaRTX0W1KTaRWHl/wEPmVSutJfswZ6ik
j+nMnmY9Z9Ks+srJvcJURWri/goL7NE2UFW85gGQQbVbzxp59UTf/aHtbgh3MDci6JTuCDUVrUoB
57S31xNGcvuKaIQdc2SmCvNobuzlHSFJauk2n1fnkSEjr8/VZlUFtC1oA8I7li2P10WmhHAliRT7
wIu9OhmTGMqX8uvBJ1gZ+8BvJb9d3t06gfZPOdpi9HU4CmO6AS3Wg0aZ2nN/EsSat968K83uRftA
xhX2Q6XLCZfZ246ca7W80VCcFdwIbKJ/0LJ1/4agPzKUGx1kDemptHbwsXlWN471R9QTLlO3SeoH
WF4yOJzJoNve6VV2xXpPCCccKiuQ4FVaPqKxbL03yQzht5DraP80vyiVi+uI7x83cI/C23X3AUB0
6wlvYK8HeY8RUvvqccNlzFYW5MMWyoEjLK1a7jY1vtZklHzDx8uWUc+r5+bRA3FZ4MjV+sQoS+rR
ZaUj1Ne0jHJKCtxkaNZ2clGNj3aiwlhtuva1DtAt7osYfNk+k5psoIBOlyh4hXa37+kHFtiUAWnv
qIdtlKWCZLJgxBbpdB1IsAmoVNFGzD4W+ZjgadieJxIICpmPrKA9Li9EJHzh9W5FOPzdUms3JFh/
bqtTNmYAky9X2iG4Jj53EI3YSoAkX5cZzYI+mF2Ctf1iQfLpzXfhasNCJ4uNBWOMxNhYFex61a4i
YxBlxJfFnuanldRjFGbXIaH8iHUK6ZTegDM2XddE6a2o4/H/S7bnBDTll3TeimoB8svycWNg4hlN
aRrkBykbNCnGCf9cZSJiUZngOR7tKasaZRILSZBCjRCfe5eHLtM5tamHvrZoQ2pnlooFZqfd39ei
o5gK1U8QZzc8zMJk+2p+X3qf99PC/pIeMB5Dcc+KhkV0dD2ppWVRAtJBfQWsX8cUNyRKKzB/QdpM
cR2ZIh/7AAnEc4//lkvRbREEa5371UboiuL/fNJqEl/loorSn8u594wP29RM/1kghi7XWBn7mpRD
xUIW4yZwsdAdmz9T1OEmPDRXtwsv3FmUhBnCEifH/vTvSoXsLE3EJ+ki6nDSVfNdErqVxg07B5zk
CJaIvlVuE9H6UBLEzBd1WMkykG9Vi8v/liqqr4/X3w5hsH/Ttja2by+MhvVa08hPnxfuRJVaq7ti
GcH15kRpFYal7YScKS1teE6twXCkAc2XHdhgJd6UVGjYnLwSUY4xD+PJsjnRuBX5kN2prmssqP/I
eU+9AeGda5AukicA3/mYJsUYsBDQMsvPQ67RMEh7eM9U0/5bESpyWSjAHso4Hm9CMMP86Uyyd5DW
OvSKg721yfwG/Dv0s3c0GtDwrhjreGCENiyA7aKTBjnRPIYJg+trHrOgFTsiPrKNNOCcUSIFnI0L
JbM/fcKt/EQJ9a9w48GFTm/TgPTzGQrWnTdgy+Y5QB0oeN1CymlghZuV/nLhOFIB6Krk96VRBATV
0ixKgytYRkS2T4Z9YbUNF9+RfZYTTB8Qb6s5b29Z41vtktXkngQyiYuJeWrEIKNIqksZgYVNyFJH
Yj8i+Rviavc6pz2rs6uGo0xEogtZdSQ1dmwk2zQzu9jx5dW4zQYgMwIntEcn4oV4piTj3EyusN8F
/r2/OyqgSVh54E5PNk/D6HlGpCAdoMqDHBLOLzhGYOD96r3rcXIVwHZXVAZsGW+nsCUBs9xMunXr
ST1d8tqyk/JAalcgFdsV01pHCAMlTqyHyzCadCY8E5v/OF87Lz0LMbQzXLYBMTEgNJukAvDeS0Y8
a6EsfuDrV6ITXp6STI/9yqTFmA1izVCsyOMsoc1PKT+TO60l1q2W/yIS1/FT+L5Q0h3N5mdDFvQY
JymOdYaBNl6YqvHrg4jqhHqYbVYikyanfVFFPVuzHxSuGn7QcCBmIwmYZi8bXp4z9HeN6hEdcEhr
V+7pTnzrgHqoLi3pWYYmlWYm8cFdyQ1fAYhaWLoBRJ0V60luEEktGoQgTg67u4qDFwiYR+MPwTO1
hv2BhpzM+jtDYOMxeG2fINMx6rVdRkp+0xdu9TsBsidVju67tLjFh4MQZn2RQzQFeEmLrt7kYIUE
JOljSiIFMTrpziC6hARDVE4eq7G0komQLah9TZbrSkxzw35bjnIo2p7pkQPXhaZU8wmrc9A1R+4J
QSxXtN2lj5jnl/xpdQhhxjjlQFL5UCbpMLeFt2H/vKOX2jKKbR6Ajr1J4c6Q/nuGg/iturgm8Ift
tsad6SKjZh80OuHBt2tbyS6Dj3EyUUSt6Fv0cgsD0rAMgYYWDH8EYJBETvif9fDBmlv7OrR9zq06
SZm6ycnQYDRGhuBa+AMBwWsp9WKaksaOW9GQWEtd17DgsClzYDHbAtRx5I3cx5Ak2pqUB5uYzxoR
xrOeVTNMfq0O6cIL375638BjzePhBxuqkUBLzs6bvfFXuWAvfy4JkNz4+gNgr/xI9+ioihWpN8B7
/1gue3YhBILlxuklyjiETD+8Q2BHWoifXtkWTz+KPt+ZP34l3WXJugSDPvZwwnG8KvDygkGtz/28
+bY06YevCoIzzhh/uyB873S6OHOkm5h99dbUucHTWY7/uI0Ah8k/ccEFbSjIJKpmv2Qth6/3hTRG
ROKdvmTs4spuChK1Ra/PWIg03zQng/vuH7VAAfVZhpXy4W/AKBiNTh6qSWc4LVJId1udrSjoT0jO
8l1lDHCiHTQa8b9Ub9LNMW5KOMavx+PiiBN5YFlk0NZxgL00faSxmyV5G7MsNr2UlJat7bCtTTLm
I/eml3i5DD56a503U51FNKwqaJbt/6/816Crci3VhJFt4/X7lwWL0Yy8YDSLYda2NvafXgScOr1u
ZLJncVprFAm576gkF2RZ06RmqzMTgmkXQ8zQiH4+ztwAG1HTRsna/FS3a5xeqzls00r6vA+9Uxs3
7mtt+7//JwiSqRm+sUf35rKzslGYmp+uzbbKHuTAFPR06zD98u0rq+HZlvkYCHiV6tSZMTD2FOZn
TaSWryPrCCkUQwLKNptK2febvrMyy9kF9v2Fk8+uZ8MWqNLNVZ15GP82ol4ru+CP5LlUo1Bg7Hhz
yE6B9n8J62/TLjpwZ/eNuBG0K48YVoQpRMcy+f8a/xQphJzB1CEYmJOpTjjzdacVUHFxKffly4+t
WvA1EEvs/3v6kSXyNF4W1nrtaprnCaxL8jsoFjx2anj8k/mahYQi9EncSo2mXrIRTnnOtxAOatnf
DYPViwqXJQ0GamDiNoXwrI0WT7/l4yciJ+PMQUxQTQHo+6Um8cMeKu+ucqvFQnJpDVdK0lRZtici
PjhFRb8dasiipWoKvG4o8I6hOWrSehAQdKtThwoDE4mlL1AGdhFatgIeTbfJaJAuAQG9yWw6cmyt
E6RMlEIf/ZgkTE5kV/s13erXXw6d+ob/jaGR10hgLKUGQbhWBBI3RYegXpSUfE+Dr6lcFtlZRfho
/3ftPWfB4igqLW78phQG3ZS9Tcy352LaqOnQlVVdTIiWIH20znwJI/05AZ4VrF3iehadlkw1Regr
x/NayEtp9RdBh5A5UrRzlgZD0H9sxxC+Cq0t3HkyYDk+kBuFcW+nuHJdO9N8/jZ0m87C4E2WRr7r
IyShLXm3IJnHjgfjikdZzm2GJJTviuVNzi95e3VTq0ETqb78HqsDsB4pq88pe2W7BudOOCgbgv0l
gRmSD7gH7vUUbOt4wxjVSHjDv/FmTVETNofmblA29OEuHTqKV7yLoproo6xIomhifbQ79l4yeh6d
B73tQmD/gb2KpcGJgO99mOIFjHyNv7wDfJtN9Al60jH+8ucdKmcSC9HRaUfurh8d5uS9zstoGfWe
vI92jO8iGT8AcQWs3LoiV7xVGlsT9Vxz7yBZ5UL7IIXQNYH2gm1CRAj8sspTq0UIAqHn74jcLFt2
vvLddG8VIip7y+a91Amtz4cSusMhJVSndvRXq9rls567hbJxnhN+CJuKz02UBn82wNnTwbJemyGa
uTQSiSmRidn0ZDidQ+0PJf6XwUeOYfdL2vEGYLnMpMu83Z7A2O5UyFf/1HoJNAuOk9yD49ZoEsJP
DSabt8ty3IRPyAf46vAQkEFVhGSzbF4yn9BUwgM+OF+6Ij8QOcg9uTCA5bKfWdrQKfEJQjswb1OJ
qa8DlGVSRFOd4UE867tr5rPkPVV6vzZFkLQZQLje72ApdrglA4IAHKRavJIsqqp4hDF5N9OyAt3G
3KnUzdnK/SjZiJCCeufplduHP3XI/6giB3e4oFIIB/w7SmrB0GFtm70t0p4NsQIsoi8lgSg/Db0+
HYMLsg9fq5b+ny0fsAi6oWh9+I7jYOajHwf0u0c/alNkM05jxXO8Tibguw8MtUN02tHJcY8VzdCk
MN4Xh1oIeUDGHRpsvVtUnIMf99nqFATLezi1ZX8KIdubBOvcm8DjSUkKm9/yh4VV+QwBKu4V1skm
dV63NmjfoMXhB5b1KGpVaUVWQBWLr3zyD4HH1GvRryMrgHcQVU71J7oXFRxUwoF2WkGzp7DGMigA
+eb9OIg+bplRiHw9ACGaJr7ipTqVWl0lVYJHl7wZULPgftwy5OAESHDgfz/hAL1alAfSo7RfvHNV
hFWuqr2qEFaQJhHjOamzhrCBt8CN3R0Nj5RmSw68CLTi3g57MYkKd8ogJ93tRlrc2PgHihZsWefG
a2umkc7pQzu9vsnD/COyQGXZRvfaPbGhy5xjC5JwEPBcR/xd1+n33VNgw96dLpjbMyl9im4Qwgh2
5lIVJdcwCflb7uNGZt7uwxFUv1iymxZuvvmQG7KF7JaCyT4jraZldrOhRmn1Ijg4QN+MmuiGx/re
TAzaMM8QEa6vfkkmk2iauMBPpmK6qwo19sVI48/aUecDx3ykL5/3CTZIld6m3R1czYpX9bbtzXZf
sJYAT2tUgwu71aoilENOo4A0qQCpEdamqhXlr+WxwRVa9OwWzAKxJTveiQ44/7G973R+WPJSYS+/
F0ehoaxX8rCoWtAeOh1Y4hQCprLr/l9wrCI0msdSsEbind77h+NEfumOTiKeBVxCcqst6x+bgKrB
v9D1Whrzdcx4tnNLme3vOYtcXLq7iToyrMZjApLUGLxbQZ///kLj6pHvLBG36jsWPVB3kS6DQVj1
MRXlgPRIW/d5wxe88TriXcA0JE0U8CBMP0Bvr9VRMzeHvb0ixyuPPuzR8vLuYjQDQ8IJpnEDvZhg
3myuC+dbi/tKPKnKbg8VBg3AZKCjRhDMFPiUn+T3M50FlvJDAAdHMsm9UQdMCeFmVXcZiV3QUC0n
gv7B7larOOwa2mjxOlpbapztgeRc1LTquH5Kjq/UIrN4ZYuQFkA1QHSt1d+OBGU/+QkiLv73oA6/
Pf7XBcxQRGcgF5poUVcbOuqna/K9+6JuPMEFV59h1HupQDgtrl/golmjptSGGNaUrlOtFLXF1R5m
YzPkHXgoRCh0cwwgp6N6R4bucb/F0Vr8H2AVuadav68j1ch8JvfSJZ+WzZYzL3yLjb74Z4txNyzh
n5MuMu3s0AOzkAcPaX0rY1gs2GflYmSTBMEvqtMGZHGzHVhGSGBUpBEDilIthNJV9xUyqW1SUk3F
/selwtzVn5uA8SrQGiHZ41/RTJmBcbT8OyTsyIblR9eZIFBWbXX4ZdbIqGxZtiHVb+V6qwN4XxZk
CJqBPKrZPzeS3GiFWt3PQGCqMB5joplN92B7tbtKXcnkDVmwqP4WUDDg5qBEtkNQ/YWJ1GhAwunN
n1YiR40slmVO3BDZgJwWQ/jaVI1Vom5+ruzGkF1xLCfuyVYFoaghKjF1s/8N+8gSZWvuNcww0Y2q
SgnB8mElzsDZTrPW6VzdR9TTmOQl+xVeBxh+SYQtimXKlnyqWh4ebc8DCEfR1zm5ccyLsmgXrc5c
JdAIa1pMlKZvx3CAD+blEehULt47CP5WezkW+Z/rt3PkTp7Ab2gwkWA3NQIsEMai5HT06f4GBEi/
FX+/nNaSgbg0k/Z9e9kTeN8eR9p/vGy4D3CEMRbka41SPsMPISoDYUTaTTSxv/r4S28JwQnD/zmk
uegfq3fA3TpijNX1el86NSdiXXkSqQYcabqDbH2OCYIe1hSvLEroPGcNre883KAHDb5hETY27VHS
JJMWdE4DJTiVYJYhSiJC+gOGBiw2xg6VDqGE58uLUPAr4YZwr6N7EjoHrJ5auRBPgD5j5f3QRQbs
pVEm7gr0qJYy0wy70qm4140M/ENXT9fErsOBczBfe5ktFgfC7yNyUDOGqEpzO7sdJr3ZTfe5Fgyh
3DkVivoseH8RwLVKgXBfHepBrCJY/FUw/lFXFTisuzmSTYAFs2wxh5J60FkQIWWPrrhVii00laNP
F4PPAC7BDV64y73Gc8Z02W822tFo9iCHj4k1tdTl5HkLYCt8lsCbpWqMg+yzcDgaC08qc/Cl27Y3
jvZ+xyXB7PE5Edy/ZhbSQX1f8M0WRi4vyN/3MVFg/2hRldQKh77tbj/NhjZMPBfUi7KzdXbxTOvH
HykMvdlDQN/eaHADrPwMuhorJuQb3LeWx4VqLE5ajI5/Zx0OZnG8eU7F6wakW5jJPOEJUvLRqw2i
GRqzgRHKIUtdXKmWuHZQpkfuX2e2uEGQ0yCHQzPByPkRvB+RjhrrYvxyQ+Kxq3z2WWapOuxV5Kd4
wl3v8Twmlr//GmnYGDN9hs4cNWw8HyYTuaJo8Pav4l7BllSoMCb+yC/n3SxPV9w5wPi3vQcGJHVO
5TDYAW7To2uVe4xAu9ydcWsQstwgetyhZz1+DM/3Pi9TLlyPO2rFA719n1gvECtOo9WBqDXsamzC
+g9H4E2jYJK69yq+NwRqilNKLuLLrmsqsnRI/mhsuOrqXEmFOyDHYW2n2N+75rTJoZcC5sLPX4Z4
AvWVF78awbIbaXJppCy1jJTJ41xW5s4MpFlZSuPXeuIW843FilWkaH9yNsgkNRgBAN/eRsJOSi9+
oCFth1Mlvqr4HFf6G1u+MuKe3SmYIb5zkjmR5FZVt7Fn0qs/kAHVP4R8fusr8l0r3ZGpWUP0G3S5
XCMltpshMVIxuZCDyYoWC1mDc8nHCUSVbzB5PkxpYDOu32w9oFQAEBUezAGI/Oih6YPleEpPmf8x
lwJlGrY+LBaPOrDGSjIJahDCLjxnGS8jFonRREHKHaGOxAjm07czbIzLi9SpIAqbsAi/d7L9BeqP
6z7Qp7R12rjcmYiuiRsCj32Z8FI6Ha+tWlKpJpnGb0ko2ERdVtX5IFLCG9+iUkP7hQomN0ffWw5j
zI2WRw74wbNp1uoCULd0q2/jq14E3bwm2pGnZtcSro9F1ZbfqPTSe+FfRAGDr19K93CnMC8/D/cW
IL/JoO8Qj0efH0H7bn0k/Nw+ixX1mBg4nqh+3ZpKbzl7SGHb/0RgnO+lnuk+f58YOC7WqwXOy9La
MtUUeKnoPSlx7rC8etW8w50KmNJBNpN618nvz6auDo+lpKQKClXEis+mS8bu9PI3kSsDMeMlVsvG
Mex7DlduzRkbUgY3/MmSJMFg1oYtm2P8rsWsl2IGokHwns0LeNZ0nveZmPUOqwue2eTiB9eRMyBb
hWUPdHEiHd6IeSAe/En15qAlGgi8IOAC96vmCRtuqwktxLVN/DVN0rj0V7PAlFIzKXSvInPqyIHl
DUl862ZhmP/nk/NqEgeVspVahGna/h1S7LQR39dliX8sLh42H01LiCroEyl7SRkKb86aqGA/ZTqj
z9tl06Nd0CgNA3g3F5/EN8muyizL4TMn1n/sQHpRmfYSW4NwmTcRy3cj2oOubmjzhzwG6ZInXNy9
ebMKgzgFX3M7ZD37zgXIgfjK6BW6m4qA5V9jKqnOZ4ddJ6TJiPNtilxeayuAr5Mi6GgbnoK6kkD2
NFJ477x1X1LucomIRYF/vBObv95eAVOKNm5MXerrBQZbNHGIxwZ7nyqo4ohaEc+zy1qQvRnet/m9
zjS4F9y0sT5TkyzMaVkJQCagg+OPbY84GgUEk44cxH8yWTp+1B5eY2eIEXMit+NTHR+94bX0CFGW
UGMCSLlaZXFhPIRQQQvoGgsnoGm5JWcqiHz39NmAO6I6qmo/zRjoHlhXQvI9MEva4IKOg8Yi9nir
/yt6oyqiQ3g+CfSeP06bA1sPOfeJhrKNUlez++5Ens1Vldvg2GQkQf+S2vaDhwcy9PJrjMngAV/Q
V8D5tAqvLPazJV3hzyKuSnUqvEC1xV9yv3Wke2furDEVJyBR7gy7h4GLc07XlA6ogEjAa5++/l+/
nCFAkP0G870dG2Z3i3lnQsU81Al73zUVBMM2MT15WWXR+kHPXpfj3ed/l8s80244b4pI5stYRnHv
N7s9z0zls90939hWNX8TN3rTBE4MuuHbZXURjSWIceXGOUrd0xUUZNf9eAUGNfRezCrFwSEEBW6S
vqOjLy6+a5ZqOIoepHa2NPqz2JSPIEBtZAx7nbvOPgwEimmNk/QmccUlb+YCEOzzO257dCg0WJxT
acxrfNKJTljF7RkW9AyO26AGHUhwUXEK52zOEw8GPRCXZKsE302YW/Ah5kMULHemzPMBUSRWPUjV
d6FVOSZ59H3hlXMQNXkmB3IcIN58QkFa7JHPsMMKsZkZnekFHrl/ptX4EIojy4ddQO37zcEQZ45P
eR8f1+4ABjpF4XU5v9b++NnapYUdXGaKGLeNgGifgeVdjkHUUo+14GWJgwCof8vMMFLHfF8/vwWD
LV/9I8I9Xlm6P2xrmUYVNGSv5EjO/HZZTKIZE8w8If0EGCrBKv6aiAwui2+cBsypYGGsOKKk6RmC
Pnd0DuA0WxrfSW6ZehREHi8oUeB6B4kVxU7cPP8VZyS/ost2Kb1RKK1JF1SQMs1hrIb/iv+OnawZ
9qV6Qm0yAtQ6EUmTYAGFBLk0112zfcEDEfCPybsOsgb/BMf2U9sjx8bRzpEZmVWr5gN5uP5o0lHX
54R0gOA48MtGyC40NfNldxSrLlNOCbQZhf+B+oxOBO7lr/NzVOVA9+CIxhJpC8k6TmtiOFXEZ0B6
tS2HKU9t0JC02dh4loauChAUmdMDGM8Y6NSoRUi4Ax3wFO9TUXhfQTpwvp4UXtcTkTfmTtpkDRWN
dJ4Flqa3j1QFuMu5bOw1QyPTFD5ymkcyTkStX8YwPWXF6yvqn++aCVdItg3RPdcz24jx1kqSuTdF
LDoGMa/OmLQjVaugZPuUOGGxVc5wjAXLn9ce7k/DWWM0qcQ/7V13lYAGKL261xGXD2DNQmTZ5x9B
RqkhLUkBzizkEu6QBJDG1J8kWTgHTbsUqG4WpLTNPSojFyUD6g1mRU8q/dDW8Lkje4fkOLHSjEdC
KHYp0OCtnU0CtZaqLprdf6rzFRhiufjyoK6UnaV7yopnizfmoYiK/toj5i4uPSIQvqdGTqVOBUQp
tiRBMI68r8wp54DMZF/BY6uDMA6MLrS29RgBlCrsBILvIhOVSLOFXMQbWM+XMaG/4fRFLm9N4vnp
TdgqKTu3BEYOvGOTDmD/TNIWBhdzxSW/hcJaSU/b+I1laDSmEgAlqqmpbUD3cRbpcKM7438pKi6z
T0TTTaBGBDmMct/xzxjQPbuMZ1mhWbZvJSKE+Uybk7UMUsyKt2vdHbaFww0nNZI9miCdl9WfeBsq
/RckId1a0KTvETS/f6shKk0hHksACVMrGxxb1Cwc7pGbtfTVKgJ0GwQhoo0B7IVuQeZk4URmZV89
XWh21UbjxbQkCtHeCxXkyK9O6FCQl8m7hECOkaA1MM2j3iY2xmni2pgvbiW7cDHBFc7WjWvS5TLs
q481sSFkIRNo/JGZEaw6bh22y9bre0zrqkn2AGicuLa5gl1i4zC8TrhqAxLAmCosyMfYXQ7FOhUh
4sQ0qrw8YUYEZ7/jwIT5gqfJtn2GJs0+In3CJjScnNlzumxXzYNgrUcQNoprAZD/Z17IxZgsYfy5
ImuuR/FXAqKd92CwsLLiVlk0rxsCf2syNdEKVt631Gg1X9X9MQhZ0tTHwvV9syFe/qi2KSdEJDVh
K28bcndGA3YbnYputUoZQMZ/0KF/XhDfiZvTPQVQP9f9rZYbFPeTl7BYu7Cevbnhd0KuWrhwGYOv
uGaTJCNlkcV4VUX4u16iRPXG2M+ZSZI96mexE4G9fn/8pm1v6wmpQj/JE8elgY624BKj8jMVNvvO
/gD/blpm1aSJ6LLCOQchQc1AhO01pER/QOi3O71Oy1KED4Gg9QIVNjxqVRlcTbE/ZYEjdUNzp2q3
n6S6ex7EjJcqvVTPAMaSZGXiXVpuYhNZQZ8P27aASp9eGH+ilGgQh0J9Ddukwm030pnp1llNAJ5A
hNJz+UjIvEe7kBudDVSvil5xlWNr44LVFN9lQXzjP8aUuIY8y5ehIkOYcFc1H+yIcNgLPh67s1X4
thKLlETLNl6e4ZaQLKIYiG13m1Q5+NYQLHbwA5qRHX14PYk5kzlrasEfL5gPqPdfkDPoXEh85d63
oJMR6o2osO9ct7Kq2LH9dN2X9sNeC8AkLOCi/74EHCcFyqRXJCIQCMYTmWuwlF8Hwq9jpSEYyq7p
d5WOUusWzCrh/dlcKBvMtdJL/bg91Z/mwkHjaze98QwI9a88bWSMlT7UylLHxNqcuq2IVj2z2puj
2q1edM62QEWxlIPFSA8wEEY439oPOR0CdpIsnDvg4NDaFFm7YHLYym7ylVOrUpUnEyc21pFKev3E
nwVqoPHNhAgs7I4r1VSdiIzOzVXTGjxEVEk6JWeELig0PaPFfwyE4jv16SBjyLxRVsT3hiQnX/1J
l56W9EC8vdtbaprE30XurVYQexBt5giKLz0cknfifZCex7Km+kr9ogjlJLozoddTiCPAnsCec4hs
AF/VITlPFa0lMXJIkoCMP0LhtyM6lq14OAgZRKCTdVAT3pC7sCmVF5z6tOhVewcHQEg4JEDl+p/D
D0oQ68nAXlK+pghlQs7vV6zTr3S/1wzFmXHdGpcziTYh+bW32TAKmfmZiHV03fsd10So11jIqdSO
RacBKr3NYp5Xs8L6hUowKLizuvbhuRVTC/UfQYYe9af1AYUi8ozbIQzQgXBgU9trlEoo9iu/65zy
86L9cQTc0c2uldiPCS7n/uS4rQXmukr/1BCUYimZ5BAdIUx2BmcbkqhI4z2frJoOTs0/A9JLk9vE
BuFRwqN0dIMebPNMmF6HLa2/44/cFy+0npwvmKh7E+nUGGzi5d/38UnnbbkaRzYZCX0AFM202+lS
6xXRrxRo8kll0zbr6ooIa8/dlrXq5aQoUN2nIy/BPWldseIUHc6SYDmXv0CKIR5uJz4WlMzr6gNM
d6gUEltn7Nh9oi5to81aUc+kBSAYhS/+bcXwCwtxHowe+2p5p6J9nWtYCMERcIXzea0XZAxvQDh8
FYBk0Sk6Yl5/ok0dGMt8u5TtXYoOylJ+IhY4YhON8T5jmCnfccFfLJQGYiaqbmjkU3pvintleGUO
Rbc+ThQ+keChZYapuDmllQJAL/yPAFJ+syum0PG8reJPM5CV5SspCKnwRNLbMa3jvyK5cJk+nAAE
HxJcfIaWay0J2I/kwXgWvJKP0DGGGHqhHJ92I6NBY7Oi7J0gIjHAh/z62dKJB4zjVE2Xuig4Mahc
Vj46Jnku1kOhrUGGqTaa+vZfiIBTM+6gLcKFqNz83P/cZvWSAb5eCiQOs54CaztSCArjUbxHO55Q
33VyQmDoBoD8bw4aGOSWkiC71D8Pl/9Yc2s9i3KRnBHi63yxBdz7S+Usxedtw8fNhlnbsfOpC9x2
5FDEKQqOCQs/8iZIWS1Ex4fkq4tXVtH/HySZTREwVpMLxmS4UfsyVvAUEIQUnIKE9uYkxc/S//Ts
nUvBvI0u8FfqMp27v9L2LAmGTxieLUVkUbxgQVoRdudXaQSgzp88e6JbYU+3WBvM/UNydYDkCHTW
1x9EGzcfbnCy9gDBnOHy8rkp9Qh7/wDiAf/q/ZC8HoO+eZV9keFCCslJNSy4CZBnAaPUk76w8CfR
npmTNYuqmDYUfM0YKjdQzi5o/sf8a8bwu3q2Be+hJVqJnF/HIS2j8y3DeKsGaOg+eUTWAQXrEn3R
8XXAQzKQrN+/ZU3pvncX0kIeUC6o0tro8RpNN76xDv01amfPnvviMUUFtXSbBIrzUqrGE5cIgpkP
x6inE6iCoDmir5Xi5yYDILmiM+s0u4zwjCMSlSMh9ZL9DfrmGa6IaojCAkgJwg41S1iPUWuGadJZ
YZjKMDK0uDIGuyPA8VAeV6RDWwCuBO1DaYKWl2e8/A9iUPZe39/ro8wKDpI2EEraWRwyfeI/9ThT
s1DelR4+8I48t2sZzXbxWGeGq6CYUigwxRLTjv1cdWzi39TjfTdmp5PF7GbcsAaTZfITwMLjpiC4
Ba7XQceZgOxUzYzcnuvhmNaXG0h1CLIqvtdDYVWF8pQ0HFykN1oxG8AMPGSj1hk7wsO7hiW4VmKL
vLY8aVIBkoTDh4k98xeyTxRcmxNG433nAVHiWJz/uG6GBa4CMccKaVi4kHZESChNakXX0SYBFcH+
7hohTC8s0WxiSDeTrmRLjM6WF6x6kWqq5qm6A2tHPPp2Ok5KcpEitKzUNkOtaaWoOLJUc10+cCfM
c4L4VgkzpyfYfAWoNJUyKge+ejPNpYA0ixTolwDA3xO7UORnvRDFtxM80ro7FljuWp0l+FquQgKM
tK6QsPETHBEFjfNXU+YhPoUxR3qQ06rjh+1Eo1FIdIQPf3H9GMT2Ov2xq3fhjT8QgsD2fcH81rY7
c6++fOkLoci67EN1E7Q8V9kZ8vUOnBsfRjJqQYCkl+966CPBIdC+s5KB/+kulcxDnZtAdCeN9UKV
epOS2+CZ64LI+C6Q2I0xyuyzkVBXT6lH440UerjjCnTnbY3T8cm5ZpfAH6q4U8tdz7ofNCKeD3V0
ThVL2uPzQfThcacfqSZ17jbzOwa/1ApeTpe0soj3U8jZTyYevxuHiQkv09FzcQmwl+pB3En+X6tK
AN9VtyImhq71157sG6XDuz25dDhTC3g7E1wMBouehfeK85dkWSeuYakvB1op5XNlTxro+muePdlS
/Hbxe3XLpe0SjGFlIJTQDyxsKzTwgQhrXQwdNiws4LMQgk241Zf9z8NIsJaBKkjElA2jaYiTgSDI
KbNf8lJ9GOq1lL6wfs2pUyT4l/CJ9viM9GdnHYO4P40qFjGNz3KdYXxh0UG1tr7qhTSIMMMygwen
0wk6i2G9GFoN0Esq1QTpWEHwySx2zwf8QlCGb6MRtj9XHGZfKbqtj2ssBUJv7Sl0/MdX//fDXqA4
+l8FSk/Q8WyzCyDn2wPl3lrJDh5b0qyPiR7dfAEAzAFmPFAL1aNgtoLXxayOQ0zMmNfqUv0pizeW
hKqHqhVfrK7/00P6Opc4uTB5DoXxcZPKSxXrDqOUhL2EQc0Yyv1fUva5k0whZ/kB5wliT2XTQQdg
1PLAQvjR0f5GDP/2O6K1H7wOuJiDZ7zrA3jg4GyjUtZZzOypXAHzBgVatvDYQfgKWJ8e83cpV+LR
OMZHub7aEMJj5FG0wTh5rqoeOV1BnJkwRzZk/pEoA3Goqgxn0UkQdhTtYE9kdAWDB8az08UsEjCO
sH4sPK+Al8SbD/09m+wuFOXS/unLeRIc8MWx6sKpAp1a3mpThpiPGczd9D5Q0KA3+dwMeMA0m57U
hQ1QRyA5sOQ3N31tS/ndlOkrdds8cKfkObzFXpmJ+PP2s5U6j4gBfYZjTanT+2OTAuWiKEp3v7rh
coeDTrvrKFtaztWBV+UbCivXGNF8WesP5Y8beSbW+uRJFobdGwToLx8gup6c/2FFPk7CoIkTW5qr
OpI2dK8LYXcNII+M+VlKAoDwk6WqQkL7RUlPIMeAxtoiCEGogB7b4ORsUVAuhXLMm2J+WMoWmUx/
XDOFtmjWjTk1AGj2H4fE+l+z09iiq1zd8fIFh4JpmARcmDepsKlo3HbKmcPKbcnBUHZFOjlgN7tn
p9IOK7Q+UikwtqQ8VJwpf5xQ9+x4ZKtqcI8GDJJYPP/nXSOvNScg6WV0e0Ax8CCZ8eFzBVfUE/z8
JpDfyrma3zR+qGsmNSgkNz8YSLlqMVjtyYlYtw20tUdqCSO46pYW3cN1aV6qZos7rqqRlnL3AEhX
EZuosSdbE4urip67V6m0YZdEsH+iF3iuVRyaJPWYc0l9BFvlXa0c6rd7zFx/V+pQGtlkTJXPGyCX
q1gSIc5umFHrFeto30hhH5ZknwipzWqa+4RXxlakiEYMo/UIrbMa5PUG4sZZsYmNfHY7nk0AIzXJ
HGzHhZP/k3pWnDL1ip8zzVaqPb8NKGu5N1u5p0tzFd55sxI1fN7g+7ULKPZCzh9z5SQLmAPBi9nH
JPmbppwhngq7HG+wUvNHaQaHg8ei0bkDRyxGSjTltgOikN5nIa6N2hzBuhsur6hm6cPoU3+AgW7z
gfVi2zufBJ18KgK0T0RvsiV0MKv/shEb6o/yyuFYARxUndG/N35cb7cgzMzKUA/13fCKCgV55JNC
apVZwK2ZFpbBlQMiSYl+1Y1Dtdm7GybxoDX8/QEE8AHt9VomZQfP0HQKW7IL2UtG/ozgV6N70DMB
yfSnb5MXw9jnKFncBWvtm/jtOW1wSu6/b0eguo19ZjSySPFsyHpzPVsFA652AzJT2VWsKTQNWxYm
iWxxsc8T9Zil/ZXyFMTptV8N4B3v4zc/+5lnFVAcn0gOcx58OtU6XnebhoXvB7w+VWfSNXdFHXKc
nIp0+U14sF9+M4g4Uw2ZlBIapu7l4+9abWVszx1wAJXublxyFeH5/K5cF2i69RX4X1iSbZ1WcNjj
KxU4W6ZJBG7r8ZJUqoT7Zq+igXfVmKcWQr+5YuyYb3wVx+FgXP8DrhFkZv4RwNICv41yhr872Bj7
fK8/a+CJSmb/9xqORWQGlPMEyk4YSUYzZPRaJhserA9TEzLMnpkUelLCcgsssoey6ylr9DcqPT+A
/oTUI8B3xPx6F2qNrnv3kEviYh5pxm7ecSg56mar9sBaqwghlRpcrS0I9Ku/z40Fn1v1Pxt2fPft
XiL0wvHDuCnMy8oYQWNod7AVl8Z5QguOOTkhhcEn4v0keTKTPBjR5OpQjA/2azmgGHmNY82E/gPE
0NUaaoiZQ/mUvlLjFctzpqIZy2uViRGD8ZdMEIxwSZsi2NqyoBxsDXTyJIRkL1x9/ozRyv16V6vG
tI0cPZOL7zOOp75C8rGtZdc7XKYG6jWLx+N15hHw2J/zkC+AHghAXySPO1kqN70eNzZ5c9C7ue6D
kqdICsfu6Pstb9BVb6oPWSfr/ja1xc0F7pGhBhk/XGAA/DFtPr14fv8qO4XfIN7cm4gBHWrT0oPK
0Lj94WzhBZu3ZnOiTMVRekRRDXXu/mgIQ4bDA7cYLlmlaNCOROI+fIlLi27Yti1TNGaeKR+QFzHP
eO5XA5AxwJgDAc47Sx5/WLf06+vPil/jNAkWsRNtdBB7xyW9rSGSSMZF5ouXsudjHuHfNmcCz2AK
7vWe7STJXf7sgEIBtKPL0dkPSCnGRdBCdADI9PGmbfxcJ2DMertTkTugU0Tg6exFGXRe+QN4IMzV
O3uHW8ferAE9C2WhacWUR/vNbTZoKDL2cM9itWuAv5MLkPgGRYflHneUpsK681u9HnUIrxEDj2aJ
VfrMnwgb5+jm0sW1igwmSu8I0e38Va7c3ARFkU6z5Zjm+pz5Eokau0T8feBE/GVjUhYDzEZKnHii
NiT8bSIpKnDF+GRLFjpqy4ISOp+sjYhnvNlxSJUwEH+PxSSU3wnEw9BIbtb5zczalPpih6XUehfC
GOtGZHa2H4GuJ8wiQZ8Hj/1IiSCkYdTnRw837SJUnHRirZzZS2jAz8MK69ZFvgoIB6Om75WBYJsA
MGIOtpqlpxF6sDm2tt0XF9Y6teWzGpxNVcm/J6MMFQeHFlWRHFROr3oM9BvXTn0r3bDTQr5ahb68
YAqqOM3KNye/BtRWU8LxCsTQ0djo0ijuGx1fUjuqHk4tg9z1lZUMqj0fGPQ0gFr7s57R96Gm5Cgp
Xzo8yYgwk8nGPRlo6Gzly2PTbnhQu7tLD1RHMRvmMM5449Bd5c2lYxA0Fh+ONsWWqhzBic9AH+in
hseHgra7FuSHyfEOqezkm5IkKOLvSM++hs/tDi9pbhDevRps8I7AKC3fOrLIM7Py9ECCV6QhPAg2
sx5gQKmeu4VStSW1DmRwI1yvNA40shiV46VYogmXt0fM1tgg/JvJDnp4D8uofQgGGQ2tt+iPJlw/
7YJ6cXFcRedS1L/HbItzlrDdtoDEQIwrgg6qA7f5gglV7zaVArWSYqAEIVWzTeCod/mqzk5x4VKc
/3XVRaJymMJ8wuyrnX/mgxN7uSzoLoO3p5Fp4gaGHSiNBATA7shoBdBSz9I54Br65kZevkn75h1V
pwh446w3/btHO57QHhOtARWz2QS/MjGs+WisijR2H5NS31q+VqYiA2RVId8ffG5eMo10+cxdNn4o
X+nC8VaAWuGVXvHWfx4IvroadBChlcF1y2T2ZyEhC/X5zliYKpziVWXt982Kx23SSD6CMrWeC2lf
epGrNZ4RFm360ArFYUB3g6L6do2jc7R+c8029E0kyE4Ohi0VhGK4D5/wKzMCLkYXdzP+5+8in+7c
kLwNtuTzcu/qtVgTNJkJlGCt99KPq6HNPnd3p9tYdWopOGARhQcuEIdndtrLMry+LGp415r9qZQS
CWry/hhs+CAMotbztsdkcyQemK8LMXZAhOWd6KfjQYiRm16TLfJ7b6OPWYStFqb+RZcr4LOA+ZvP
6TxvltV7LinV0RhIEEHozKXjb/O6HnfbCm99Nsjjio5uiGdDGxj793tOkPRVg4iDL9uNJX4QAEb4
yCwh49FE7J48e5rOAxyDhjJ7hA6tjyfFFz4GZP3caU8Jo4n7H9cKKJRHPWuWfWLkKRFDMLlOsoDX
uPmrFnz6Tz3nctYgAirxHuh9q+J7JGjy8v1YpnE7DihR3rIDaUzZyn42XZPMPH/ohV1Lc6GZBgTn
xYf2dInJ45f3f4Uj5bZ1/yXXXVL8yDct1Qo9J6ucIWqlaw7MKXhBBmMu6gakJXorWfXnc3MvW+BR
FD5CAfpGL/Ufr7/AWmMsaFNRZt5BhyOwzs41JSs24q4YdjR0RSJsX4MU4NswtHAmqkJGzJtIWOtZ
6q9BOVxge0oc4qR72EnGlKXf0Uwhbrl/w2xBkcLrIQ3wbLicvfGeqVbdOw08zD+2wIDFwaSG3iCu
HbAE5okNNXPWgt33aHId41fdRDBDCbBV0hE0y79CRAST5zMiGqyAQVuFtLv4NON3Oh9xj3fneJko
Z8b2wA5ZVpjHOjGpsAsVvMlST4EWzXioqr6JrFmZ3hJhjrouDHb1NgBBTScmW8BYXl/+xhU1umH0
SNG2JMjjQTxKklrWw90uwB0yDPZGfUn+73de91wm5m3bRD5d11Q7NgaHguMXagbD6/aWkimHQmxx
kqn7sbUUosyDtQjUUv4OZkRolV5qJgRoCZidttAgXLk7S/P+9w8u6KV5UA7ler21LDfJHHZ2U8qg
MMiOJ4kskBSATq7FINzKNlle5EEujpauH17qi3RGUCIFodge2EZ0yVU4K7CGQK+Owh6Km/lTzbRN
0YWKlWmPH3IMxR+DD8Mm0Id/CrEIIESjCnGxEw+kd0lqK3hpSaE208zAb6L65LuywvDO1KwLljMZ
f/JcyRFwCMTHBb8tt7N6REQGvIvahWmK4buYTJ6PJhzJstVrQn1K7LpusiVz/Kivr253WkiqO6dv
EEYBhPMNhg3lnDvpsMKFDE/r443Pbk2R85zq6LSnzUo6SjNHQgI4/ae32nubrsQB5yhvR2vUinmp
C6AS0WcZr3Hfea3YCbiLPoCPv6Q8jIJqjU6K23VVyzDLwTyeI4vbtk6Iu04XR/WARviIydy79b+8
c+Hln9SIhZNeOuTXoD08hpJ2rJ2VRRnM3Hq7Maazl23QjckSFDiyroZa16ucQYguSW/J7EsavNJC
m/P1etZLgpgvzxxsM+NBfb67P6ezXxtox7STq34lwwwyQRS+3PQew7xWaQx8ZiX5PwKQfcY2S3NG
jucVUiQFSNSOXUNSkwvXkDLsYN6jCgd6jhxzbHMF/DKRpVcuSM48fLQtWHzTNoC0embEVvnTiXTZ
w141P64RSdhwpHV4cAPmiIUfAlfuqpte/ULQiq46K+8QxBx0MuzeAEjiUhVoxxvIuE0N3N7HMgWd
6VggfejKdtAz/qOmvM/sXpHuq2FWD96Qrvru+My36X4QXtGDfDvbNGaQVtrHzHhInyM2aqia+oTn
KS7luJLOmLqgpbniq7Rnp64y2uZyYRGj+MSmc8D/Vb/4WJ2XtDNn0Q5usg9zBwIyQ0ay7GOgJC0f
+huEF4pVtQYjQrWmbMLjtXJ63pTEuKA/XCdcaIIB3ILCzuBCqoWSj/A3Fl2841b8UvaScK8qVbcN
pO/Xfnrl4GM1J9tACjdN7lca9V9OKNcxsta54HrHZXJ+cI085fTieh1muMfI3j4V+jrWUe/W3BjP
2zl4idXDP7z33ph4P7YsQcR4jmRIHciND+v4e+u32ZQIHR2YBaFJAah0BGmWzCGE8fUlUjwUdbVd
V8ouNruj+Hv9K91ez1EkqsIubxuIyCsuy7yq8KWGliyaqQwDdT1hz7W0RoLg4k8kM3wY/KLEpcvT
/bwO2nijr3n6BXWWwF/EwkeJImBmnSf+Znwqsm5Cn2wvhF2rIgC+APkov+74aRmcvfY2YPrNDemD
pFYUS1W/GIv8PU6Uz7QvQpFgindehCPd3XHZgfiPmxPj7kLC1ADY4S+HXbsycapJAlObl7BykrVK
+oYRQ5BGalee7IrTADiontAehX5C8fJCdnnKofirKFG9dgT7UZfGlFzBeRRYnfh6453GjFRpTtYM
RxuffsbysjgAXQhyurStxEderkOBXEgMavOyWb2Qagl0dbQY715/iYPLjqQhlv+6HxIHXIWaTnk9
agJ2ziJiGqoQEuafrZrmSPRwe2ciIqjk8s/eyqpwFLLYFn3MMghaTsMS6z5TkyEFb/sYo1gcs3Eo
C4AG3RikKKzabiWmvigL6QLa2E29yT25IY1b314rmuSa2NcwNxWjrgmOasUaUTsmLMz85Wninjkc
4Kt+QbVGYthjyPZBQbMyyLVC7k4/UkcJqnNRFBn/ZCvXtn2F/OYNo0G2Q8A0Q58iKFph35YIG/WS
nTWBl6QB80GsfwcHEhGo6e+vLZvuS4blZAuIcoXnjn5dnJ2OhOqt3LokOIropTPkN8x5h2PXDSXr
VlRUFcwEw/PAObizt2mOs90EiJtOGoNWqFqgNRyYlyKEWt2aawV4WgrU7vMW/nBNBY1BrAtO0/Bl
ymKj/U4bKIKcPdjvhpuitrwzwdM2/uSP7hEVsFZ+WB1qKTJ3mxJj2WvM2xfUhk9RGwHDHzuAyhTt
tX5EaQQ0MeBOR88V3fV/h90qIzT0vCibOZeNXLdfMYbyyKNX1uqz+DiX21L6yURw4C4fQH4XXATN
gMHgE3dBg9asxC3FYlLDMuMLUL9VsNiNvC3k7YNS0xTjY7kSzjUKblOSGjY7TG3XSdcQTTghtJAz
t+ryXV2KDzXDBVFleiBg41EbJw/l9TI/SvBnBxcfiuTLgnjH2Qsu8FggCxxuDfUUMM0PnMwn+NYF
wu7Prnp8o9hppAXuYH5EhfXkRZGi+TSSC+L5I4cEEZE+Z/Gwby0waczkRrYS/w5iZ5zhG/YAhK3J
lYjkot1tO2p6U+eYLU/u3w3KRTpknLKUS84j0H1FU4wU7OVFLov5Uido2l9PnTae6PHQrcmDLLSQ
42iLHcC/NIiRxMbzIMU3nxTVjOaY+rEGJ2X1U6Fbj3KiYd6l+WdnOSSRefsEYNlt6PiMDpzBcq/u
4qlKrQ4WyK+VthXD3Gmb/aWv7BB98hYNNI5+kF1fpjZFsSzKnyVLrILe/cPQJh8dhEYq7/LEH+6N
yI5Q89eXkqdpIgK5h1P6qs+weHOovmnZ2J+6E1rPsZa67CwZxTr7NZtzN94oimaiXaaR0tCPLdF+
VDONruT+QjdENy3IfVblsxauME/bgIgdpVjDNUTGXTX+hqUKt1b5fnycsDQ48J/93XfOYsZsg2ix
OKaEP9lhMgJR8iiBp6dImqQ/E13MIz1XcLZo12ytED27DO0Vko/RkV1PoZUfyfBJE465xknsZO69
jgpgt8YBYsF6MfWpnp3DumommccDrlsEa9CQRhu6EJB8zSapGSqmjgNs4Raiu/ATxBf8/suuHxUs
uij5nL6UC0sXotDK02f+i41J6qRbONdbL3j6/oMmce7iDgv3cH0YWPXL7oOcsBEJ73HFdBpTaF6V
nFbQds/ONnW54NdHRSoA4Ez76pCz5Hiu6gw5PTm/g+vw0DVqQUbQSxTsrTTvPcV+Q50K83bU4UDu
H2t257zRqaXTb5Hj8X3nuBVxaTiLo0rVZlWx4/5irZnhk0t0Yj4axvUD7DFawvKZHyThz8/MzUaa
sWPqeqewgiQDkoF6u43eJ9SrV13gQvASMXRezm4h/PX1T4o+rKbJL0ryCiFSpIlx5N/yikz3NSs9
dkJkWr62L7FsYFrdLprHdEm2+IQagHxzdVYSmr3WMH5Q4RBH2/Y8lFKbz1cmYiBfI0GGEtyQPK8R
Yg6d3zxbBVq5chyH4hCidRNKQMMoXxW9oRle/rPoMNPrDGfor9cOT6iMPOKjSBBcsy+as/aq6KCa
pV+36MJS7hlli9o26KQArw8JkMXj9wWcrM2hbCfAOxLlsQ2LqZZQZwItA/zeoKjDo/jIhhVbgOMX
itlg2xzDv1s5VuR9PHY1nrBUS1sslUrqROVztXU1a8521oa31u3WNgxJYL6UZR6EmtA1CAd8b+Au
lxerEU86Gq4bDINAxfyp9fbmTMd9nZwmbomcrg8uuyYQIU7jKlrdpF/FBjSZkrUDhHBCy7lvqEUm
Hlive01NvNdprQPesmfYEjlUiRzRs3A25vTwxyKNFoTfwg4K4Q9Me6MaqfJneav7Jyu/u3qBDtaD
7vQqdk88B1dVeQ7ncSyL8hDEwtujNsZ5VSB0GW4H+2JoVn27f9+LmxknJYIRRaNw9ONMzyvqkfXJ
MTyeumsnlaCnBZx92y76NDtK1dr8/lm/H+uTxYOezn9zAK94gDKwVta1mPrmG808heU2cL6mZDTK
FGzGrHoPDImLfjTKhIdb9VNZHdngeZS+q53ZiCDwJJIGqtkvlAFh+JS53aRwztVWLy31RI8SaBki
JiCNmwrRikXZrriVteJxUAhEx0vYvkCnc8+ZhPnieV1CXvG9N1r4xCzaQRfiTDw+/ZRN3jzOF8QO
KyQdQeSGQ/GPKQousY10QUK0b7GORRRx2tutexm1YGvr9x9RYklyZmiIiZV3bAPV7xUQO5flLqhr
siUorILPxTx7oYZZsbItC9pc/cyoZJn69gOPuN8p9zFlXpFLJHDn1dzA2+YdXUclwylGROTq1DX7
7xgief/Cl+qFAju8GjJb+5ErGFgRcUxJcnn9bZPSzHVD9mlUmtkEBKGjwPIMUr3JsAQscDG6bM0f
U2U3c/Ke8VaPvqDDtbQpECGq/0bcqhsFXm08KN1UZlAybboEFXAGJ5bk4IkwHOi9BDJY6IfiUuzB
97NSNzIxOTZPyJLu4aDgSI/op3j5mIKKhx7OovGZrQDcpAYFLj+5J+X90/dEmLVfKRMCSaAYHX5U
uWgMhddJr4Aes3Za/7SrZh5dODRb6uSLYj29W72Q3Zp7kPkeiTnMQyzBPSwHVKFtt0+fcN4lb0zG
WuSLocFObpT/6MJJ55Y8IqhTQmylypm3EeeyCQ+/ddQc5eraNH+fsd+nQ9KWIcT+ohRwP3HXWYuJ
q3EvCpyGTN4XBmmFJw7jIdgWLQpK3IBw7+1GZgicZeLollmdZPp7pfBKFOm3xikNBTwucGCXR6ph
6gNrQEV7UwcMpD+4iNt629W7zWGNx1A764rkATzWHtTTURQrb+CB4jJ89hDzsWLue8h0/+aFFJed
BxAQRGExCbnAMtayifuagPqc6bjAxupKM90WMwKumG/7GV9HfKQdk/aRdq6xoHcRZcRHaUS+Fsvh
8ljs0jw8xwQFncPk7IjabjNQnJp6vgHxl0sbiRsVfu3U6oABrA/1MqhrTNlUSuxzPFrDMLIUQvNv
h+S7faGcL/sWp2cPvuAArTfthMUoWM+EQLKMLenBXZMXmfMj2nkddlA30UPIn5K5siBOs/HPLoGT
emUvPawBNCxbOYtNTyMNGh22vfcp0o+A5dvIBA73eiv8kXihY7CxOGA3yvWeoSmj5tdPl3xxjxt2
kEVW5BMlSFt885Ph3LJEcSXjistpALXM8MRwUacrLAuiZ7sWxNL9oznd5aLbKAJOjVIG79bagniE
JPjjVNsyQKgjfVixdYzEyF6V+gPfy9Pn3O1eey5uYX6qPCYoqyzh+37j2lPsjjKt2kuAh/dBbTPv
Cgys7cX1MHCIJy3EoSa7/EVQz1uEnP4w7SWtjZWIktg2kxYljJDyIisLSKIv7/Y+ITPYalhhz8tR
bThGatySRQCWRugHxQHtVEojCoJuomxq0Hu5dY6prQSAzr02hVJ4Sa6YhlC9XxS4Ksa0lBIiPloH
5gj9aw0Z13cKVJpqawth67ESnPfFULRLzxdv3OQJby3ouyboD+dUJVCLjOAyLV494vV1DpSOvuG5
eI3YRvTluXYwX32hDZq7Yr98Q9Y+QmiRMJW5acRBwGlMNz0Qc8vDkQFYgQe2TXXz6PvVa7PQFr80
XNqizkOBkDLqtQqsPfGJcFrvkUFmZOi2KRKssbH4tFGMRhEmFcBVh4uy6iCDZf2tCELLTHAKJf/n
wHcPhQhMyW0D8xvMQaYG4F5dpu15P9duJ+pg3UiJs/p4Xep8xJ+c1kpITXFRwoOZM5NRu4ule358
7TNt5uTKcvjQP8mLc1zMUz86tFKhJ/grYp5BvVUUQr6SYXVOc1U8sL/sMfBAGJWAJmvzD5KxCN6X
52LRB97WYyy7wKaw4zh4yFYf2EHcNwE0ZiyBM5vzi6cZ14RNHoktv0GURR4Jl2dDBTynK3OSAv+J
YZTMuQFX5nlHyrg7py7WvoT7fqii/q1gFV1bmHP5f4R+PhzOgjOL12vOU2ZFZ+admhzSsPso8GId
Oco/R3AXvZ7XhscXjB+QbagQFpEzEFvC3PjCRd2iJuN8ldkVnQTSACjW6EnSRfZ4u+7H6Uuuf4aO
PZWJw9A0hA74T4sHB2LGSvjQWLQQ7OtKpEQNvyQ1+SbuF4AFLEBh8iL5MgK58li7QQBTgKGoMMIN
MA8u5plDaAxeFICAq1SWYiyyVqz8hyH/ly8/YVU0WM4efrWNpe/39Xxzdpl67dxtcSJHiLTgnaTp
dxgDA8nBqZaWv/zniKZHTmmEIAWYlftTKcZaSvbrdf6dWUtUFc4d/PMrn6+4RmLVwLAt05FcWNeu
xRE3bk+d1M/anPBp5+dH+UtnZMvvVakWZGKT5elKv0E9PKhLkL81jSwYgrCtGa+jAmyQin5ZYd7K
r3682+faIKHLmeJrSlblVW5W4GKRJsrEn6NzKXIZVJHMGpS+FColU7r4GeuDzHydSvEGtiAwjfsm
wp9m3+/xWYJwK+ayERpbJv7MpzbeCPusFh7jvGHf4G2QaqClTDpubsVVzgQkFuNeDqR/oya0xROg
q4CQ9Gx4he3gAZHz4iEtJrv11VTGkA0vcFBwfm7+iYv9BN1JRIeuUbwM9OSsjvZ7eaxYgWAIAHGT
lqbjALWIor1nWvNGgmXiaHHm4L/Q9O2IX9IUnyAQ9OvPZXRH99IBi4TAt0+8kL60HMmNgaxa7XZD
bhC2O5DAdAQyXBfbk4YqOhNXMRwoMu7hWzSZuD6el5KW4R63ZVo11D5jb6kd1ji5+Pz+8Bosigof
GYCfrOrcm36nIdYkxzHz0n+KDSku783TrRivi24eDWIwtIoHCBsHU7WyMzhIUJR7QEbJ9zTsXmI3
FH7v9kGamTTDc/vuQopTy6mjnR0HO3YgbW34e5HgaItWYgjSPjR3QCaDpz33Z4nrn8fZGoAtucHF
STwBZpzwdiJp3zaOix7bsBc4JXx7xmDE56jIPAJTXS6l/yNxVDwOVqEV/8SDOMh2tMcMc6bGZTG4
kE7JR2bYX9zyqaa2S4D4wd+q9M2wQjPwozniQuorO1+/OnAyg+ZNyPQwZBNrZvu6bt2BlOWh4lK8
Z4dMhCJ2/hln6rg97n9dIJ3/KIiTiME+Ee0SxdYnX2whlyIkPOB/hwsWtt9bUy0caDUWgC/qSm8q
dYORJ3H2ITmnwxu+VKtPjT/xebyXuf3tEWIiPZKCC5emaXX3zeXDcqahfM8QKmx25w1usvbMZBLV
dIKNFeyKosffc+duWOcfZ67a3Y9qvspsS1JlCMh8rXDYfqOE8wGHP5ubuo3ipWviU5P5ehD1gvMc
k1Joa4U4EHHRl5VeuWyjmiAQI3+9DYnqMJRBOb9sOfXFov62gllIqVCVdabZQ6rFmSS7O+vA9TSU
noYJ0WiuNB4Xc1TSc0tiXF1GlKx8HSJRVvO4o0FjaiKR86XMmPS43W7Ymv0nQlGA7+J4b8oPDik0
7g5O5hzlZBve4D9B/oyt9s7MNKRU5eUKDiI/4Jv+Hw70pp2Wmc9chyTlFb9CreyEkdLxSn5AsFLp
YgebovHHFLEqwQPcK+BYDMQIjJuo6pRllhe0rESj0zegUjv7kXmKO6F7J8Iap2ktjDy2aJplVmBd
5JN3qiXyTAUYszX7wsBueG8FQQ76WEPAVcZbsPnjtMYcIjd3T2qE5vPNj4LEb31h0/FrtN57zl2q
i4gi7DMmxejGqLWa7R0kZGJbnHxj/YzTwMi6NNuMl+Hs9Qu1V0IlTGq7kBFc6t48q1UpBbMHZocx
R6HZM+Xmy8MZ7wHzuKuI/5XyR3S8vuS7mJFKlz0ObJ9GOLq/kBZcX3KVmung5VZ24h8hU+YXy5GL
pNmzG1jhpKm6At5nNQRfnoJjdn7W0ofYiOvISKlHwmDE6aJq0ydQ7ZqkOXGxS/By2Tkg9dTe1dPs
AXv/gEgAzF9nMh/y8+Ly3BYRJt/Fa1G9Eza7fZOc6Ui3MB3GJsKwextrlJlTNSl8jQr+tcwr2ZxX
nW9e663Rnzsn77lhFf00ws0N1jgFhy2H6ElUCKLNo3P1zH01kEonJiZbgapE5QTjP11wCwOMglai
h34ZSrBY9zybgd3sa38qxRVtpzmOZWuMNaMimm7PRR8+Iitk+bIvSfsxw6DIPkCsygNnHPJI1rza
Z0fOw4ehGcYX+0R7KoewZ9LeWpCz+mF3WR3MXFSx52FO7ASODFa9EX9LQqcSCIuP7DSJcGyDu1gC
EI/U7VrFd8Dd+US8e80dVnOaTWMXJDdMFeyZ5JHpG0/+IwD3zGiy2e+4sjHTujqr6Tf5PAm67ytr
pbf19G4MtRnx4fKWtWTLsCYYr1qOodrPGgSxWFQkmfAwMXOib1VAxEUlkzGPh/8G0z9GXmXmDo1O
vxkgJySTZzi3lbi00kayP5fLjX2apM8GBnlbxaiSlxrC6SF8cS445Geow/rKQWXfLRoOXTKBOCBj
qKj9yNkISdvwLglqbq+ekN3qHKFY5jFJmnhSlkiUY9BSAtq3jJ69BxA8lU8+LVs7H1lPGzbBCmPw
oot8ydnMNPqE4eXzP61Ig7ERykSk3PlbZaQCnku2V8PomeL+CkWXVhXhnScJGAw7UZQkG6lhZGaZ
HxkVDzMx1VkEEnlqpntbzXpF+BsUZA6xcsjOY2evCzY+anMR7dhfH7cKkGLiwJ0pmhrMUtaw/Ei7
+1QcY9zOzCfgctZ/fsDzYuIJHVVRJcWTQF/QbEPhoZFM7NdORTNCiG0R0BmyJO8YUtRXLuSxrsnB
EJdANpgcpDSxbFMEDlUDIWQnasM/hz5i4ZtLpkn5TVupv1CxFsSmHGCXYQmnlh3UlCDwTVWPSSPg
T9JU8LJ4b433B6Co3k7kBsCcx6Y5uPVqhpGZ2WTiCO7ztD+8Fr9Sjuw1tXNiRyRtd9PU9UvIAZdX
kTr2yoEz0k+puypJ2D7e2HOf7fxEfbNejeg1XlkI4mVAkPLDfQrwCB4DOzPlSoygjlhnJnRvm3Fb
EJr6ywTocYcuE190qrDSYG5VWqcFhh+7iI4zlYO3yEJ+sTahlmR1Y5+f0tFF1f7HQ9WBmbA2k19R
t6jBkv6MjXMw/pCMdqX3wlMEkCNAD7jfET99i1OENfdMm36GGH7faln7EX0LBVndkX+/tBRLJYJc
24S/LMVe4Gkuw0aEtI9xqXzXcXbEzQJoVKHL8ULEiuJYIo0SIXBNG4m9SqenxMjCax3wA3+TsUUO
SuOUaQufYpzKUFupqu4eu/dHtob+U3zzzD4lVVDIBbFmrTKOcLFXdKv0E79g5LrBL3eWsy4vkxB1
2f7hBrTkboRtt3ZeiTPFTj4ErkbLQ9wkVtFIHZe9UBxzjMtLfJVGvpa2OxO61FfY4FXcE7nr9NmY
TQtISCKKd4P/mVMTUrX9/ceH2uDSiLWlEz5Mt38iFmEYHI6v85/3FlN4qgpWJrMD+otl09nXagYV
ifwMZpyXceTkPdP2rR8hFsoFOPlg+88WH3E658HKpNp8O28GhdqeL1ziIg/sLa6XGjByHY0OE5Ce
/MRaDH9LuyHOtIRV8OmNN+hOC2izSTlEWSV7LOUT/kob+4uC8IpdHWexWYhmSHW3P7ZI99PMAJyE
+BuqAQ9bTlHhTSmoWq/K3pJ5YSzbZltfCjTfRyEtTWw4zzjJfK0656pz0LIJbQFVqXs/4qLZOsLK
/lDAJmguqAMGUzhg+eZ8ameU+hfW9NCPAHTB9Y8Lw5SyxEiX/ElaeJiQVdslipe1uplUPc2hN8lj
qFuAKohzQAPUftNLEK2UetzYFZzcYKpkdWPf4sSNFx3Aa69b5Qz7KrofAmbgqkPKhYJNZfGIDbQh
dQZ9draVxkhd/xXP+E8A+hNdwTpihOO7IFxBp1ZfXZseYdzFwnXwger9ZoDJ3JA8FjuW1bvCAKJL
Ef7PdW//LsB71f4ide4kSqk8H5Sm19g0QwHliOYJgToSiLfnT1rqeW450G+x6NdzyGbY59aylN01
91jr6I44uZuO6JQqf2b9+n1VqZc6Rpbf2dH58S5JZkE/OsAc9hhEW5EWPZdwS4svzJ60aiwn2uLo
RHHUg19gWkCQtaGGsqy8SFvaDRxPjNwRjvnt/uB0N9zUVbkPwICjgmK5tHpi67e6ZvVwjPdDas28
j2zortpeDdGvinKndAAgTPpiJg0cWpB9jzJN4r6QiOrO5Q6rqAQc93XQmFfkY1LAV6SRVuleXBFi
VOSi4ASbuKE0F2qmuJ9RlIWaHSKd/BNd9TpqvYc7tkkupKKwjbQoFfuzbiDPRkOkqjD6b+rCI+rv
OZKBo+UWDdfJ/UAuGcEW5N49/oTP+XPZ9adi1Wje2QOpiyA4erzp6mQT/G8UHEVLWZGTnLYIGpzp
seFvAHeC7gx0LhosO1WaflYHvbzt44al70akvmRWhddsgdnwnVzF3E+mlZT8YjNdAdpjTSCC7SoT
+uQ1i/p20+0Ev9rTHdbjB2wEEQeYSof1XRq/bRoKyT8Y6ysZ1Xr1BXjWLXSZT4ivHiAgf7nZMolB
yCbzuzSqQdIY7iN0nJDIWn0Y/hmijmHz68b3jrz/josvRKBcITjBXabRK9amV/duQ+9Gm/TYmhkV
SywNQcoNKc4VWYvYuRtVjhwJ0qVCKvQjauX+kAIpnwnAXa1m6fY8mvB+e9SG7vU7iCniQRoWjlF5
+hg5GF3EoBAlCZFZCySulTD1i73JR94sIoIsWlCdVRJjnxq38zmDJPrw0OMYWPD9C6jEBgvl4b6d
00RoNpd63pSDk+P2hXQjbYdxUIsX6sXNCaTPVozgf0QA5DbmT6dLaGqG87AyHcyQo5aSVmbjS07d
ZGWQGLL5rRO1wah4kWuGvcgjN87YnJHdmjnINQ8EOSBbxwRFM80CA2o1+i002buFZ8+jROlRMxrs
xfZP+vqj2S7NLN4u0QIVj4BNhJNayvcoCQRUBMuxtlc00jaTF67tqyoRNb/TKOlBnVy8e0IbsBDP
j0RWmrGOw+93+Il0dcMq1XTqlrnsKdQCgahD9E19B4Hz6Gh0kChe5FfsajdfZQ43DxRxRi4G3lA9
ZpJ+yArnCYAh2LqN0Q8H/bsiuMw2sNUVsb0aRI4XRmBQIUZsqFkYEwwCHtnTd8QVytNj7w280XwA
IePVr1TCxlFTGwuPYMfkuQh3nC4z1oHxC3mPGeylfgEvcKaUMvYN7Lnk1tebVBS1DW0YGoLb6CcE
UeSPdJBrfpkPj3RspVSwp+kvBSxxrBvnxytPwMgz6Wmag7lIcYSGXi8M5HO/+AdkVs0J3Pln9/Iv
3XsJGfkZZKhEc0wLdLds9hcZffN6TckYQV5I9diDc2mZsNhqYwQvqaZDaVbTJ6uQ+nh9oFIPS/y9
oUDdUk6/Me3K6YILy5wUzGr5q8gDs2vXRIiECoFb9xLcG2ORL9KS0UVhTaeDkhFHfktwpawSBP3X
bwZf0aMhe4AtVK9C1+hEylKQbjyFf+6xIKO8/j9npD/Y/jNUux2ANOuzamj+vaURL0E2PXxe7rb+
oICevfvT1tpW4FudkefHRlMCWO090OvkRk3GuvilQDF+5oU8rRxepNkjY079RDX0wTdCqNlFRt0K
3ihq2c8paeL8Pz4xpAvNPJR8mcaypMgPZwic47IkXbwXIcalQqlu2R6RazxZ9KbJItV5HHe1nfNb
V+NZqScxQoqXMAR3Gh3US0frsQKELKu58+ztCGH5zpL8IzCS5YxbrVAIGMNszwzFKwk08Y97Qr6l
249/Q64AdcWa27x9ES3aBadTeQ2YltJzd7qbEE6EhADNa8KcRAxnKKxBPbWo9+3xA6+ojh5oXcl/
+1kmBN2XPPTJn13PLdq0WOGaajduZw2iDa+K4n03QmQEUy6OAA87N6luOD3JANTWBnbmzub/5sn8
xhdbGhTyHTRkMWc/Ur71MAW/d5gs+FYlkc2+ZSP+4d93A8/wu5R5HPjP/YsOgCl9ang45yyeuTDu
XAzLVWaZ52LQjt32qi/acS8TOTOJzdgp28VsIpN7W8suri0U962rOzsyD3eAfDF4gWBgYbGrit/e
WJzJb5Lh0TBEH5aXOZkix1r+wDVRJNjSOBmf4Gyv5JQPwclQkaqW55tWKtjWtbbnV8YEkylZqiBn
M2WMqMs8jmIi22niNBrezVDOh9csUtI3fIPsFB99qZVnpDMcmctUJZ2LnyJ6cwj5Mxh1o7pGY2Mq
G7wE5FfxUJgN+4djneA5TrWxKCto0xHk7NF9h1XV4Lub0VuWhrl/41qdPY23n69lS+LpSb90rZk8
u7hcFBNUK5ye+jtTkoyADuy6ztgKg+l7RE8Rqftb2h4C4OjPhGaRms4X3tcAzqN5YVo0WNByGW0i
t2o/jWjJLhka/mOIH0yWu+1hjL4QWwp+E1IjeRbxrAHd8IkQAPVp//oV9gTD1TkiiMSoVLDHeR45
jHqjsUDad/Imawt6ikLFFhXfSZYoV0KrPHo4XHCK4uNE148buwyKilzKKeaCTlhPur5tA2BabDA0
hK7MilzEGrXtbH7ymb3d9OHCOP+PjiEjdOk4yPVxMsuM0orayYZN1WpixDhktCKZiUtf1CL3aFDo
93ioPLFluXvaJm9I3Yens+7W+OD/bNbbwBx4OYCc8tBw30ZUzBwQxNIoRdRQc8jOTsCQYtZn9bUk
lTjZX+OAyvRLnI50yyE7FM8SfYD+77ifNz1IyYaXtptcrVdcdt2QaDzYzuQY/KM0G6FdKgBOpdHa
kXCk9i6mfQb1B7M8eMXi5qI0GMvyRsUTW0Xu3c2wfHR0Bzv5+AmL0pUvY0KWd4nDcb87fqLFIBle
nfuB8bgZgTtD7m30uB/wRQcdoulSmXqD6sixTg/VPUotNIVtt7/ToesCPZMsP9OI78byz2KDqSoj
72DPE3fAMJ+ESGdQmabzA2eY8SKj/ql1Sh6ldy9T5RCRY1sL+jPVA6ri4irowAfwyX4k582Z4x81
jRlQSyKX8pg/lAfw80MsdPM/nJik2qBWXFkyBYy/aRhInpdsNdJ0B58UPFYKMQTyLnwzBVHA9Xr9
YrZr7+L+CQlDp1famrUZ++qW+cVHlQZakzMwHjSUciNdMQM80g9INyuoxnVOkrV7PVK1zeqkuJQR
tQTYtsJI6Jb0ijxKpBRg0rbgrKCZjSGxXwhBVt3nVUIm/AtrC/iwNBAd6/ifu8t7P0+d5g1ao9jB
q2RJ5Gvqtfnokpfy5aw45KqU8z3DFKIc6L4IsgbvSjGpZajgfwl3nxSt6B4+2qe3jVEnBA365vwo
VLvGjYS1wzl8/WQpZiXubi/8+IxpSMz2yADFnEnN8aMr4e2EOFna/6+s+5PpfbpfzbwhvvFm9C+S
NkbD9zbrZeAHnkqA8wXB7+52yxrF10nZ7Ya/jAHD6QsCm+fyYkD46Fu+Wkuvk87DvknRfNThKgih
ekGRBDXNl7QgA2hxB6fTOgr7fpSTjuG+vJvdqlkYz33g7QDu854gYrfYyPXFFLL2yI51tbPSegwC
ydpe3CS6tSHiyhWmhpIbJwPfqt/Bxglb7j0sCEOgmIPV2WbwCCVRTUG9vHYX0hp7XP6RT/oxxXfy
e30AA8weMojciAIAiEehVyqskv47gfar7NV3pyq0WBfZB1JvEb9gnVXcJAgowqDICdMAj3mCfs+8
GtWLVOb3LzKe8j4+MeCjxYOdZhp/FvsMtp4J4KvvxPrDBz4tiNrlnNX9YDfbWzkJ21OHecZbtzIF
pSfRcgv0LGb/Kq+mbjOyWWaj9VDZr5YM/byUBgevaug7N1ZHKV5EV+QIO52cAcfNpM5gjZ1Lac8Z
7WLD1c/2vDVVNnoeXC/N/C+ARB53F+FkFAW44+s2X8U9YvwY5NEAd5+7vgldz2l375OzxPLA5bwy
UhVcA9C1Nv8KMDiItOORtAmx4nOvAwHLz8A2tuhRf+H24xc6zm5Zyf/E+422lFBG1LVXzoK7yaGX
nFl7PeNF4aHwOqWtzSPOfcY69Otd6pDBHuuteX6iNdkG268jTZqOzTTSTdxinapqe0HfaMaTzVKJ
n8PUsZA/s/SQdzRAMuBYif2ElAF6EKIwd6FWXDSTGQV+JW27/FErbrK37rbVD9JzP3JH7sW6z/wZ
dgWtuqhaCCbJicUOArrtjRAvVniGB4WSFk+JGirFBkIeUB05EElIw1U0DYw5vDNibbXI+4rVIAQz
DoTeDnnfjSNtrJFFpKrig+mczIuFXfyhBnla15tHDJBE9Jlxpurrkc6Wg70Z9r3pDOV97u1bmZVO
Mu3IneZEENk+jrbU5YsoRVLhvR30i8ssrQmC/Q3o0gQSFtkXvEqgRdcH2myaprjYGHjF4rjKmu2Y
TU1dxrkdtKyHYauvIe7PnMHvWXoDoG5t4fYh91jpCXJJnO2UCZ6meMyxRoasQ+tzbrzVJZr/plgU
fF7dclSb2ad2Ykv/d24UNwpaVLSiFrmw6FbGQs5nOasRguEV+U3It7Sweo3FI8cl+WZ//bfglFmW
AdVy7176MZRHkuPwMfgl9a9z6rZjYYllzS5AMDrbY/7z64q9F5Q+vNxhpbKY5CDre8z8s5nT0JgG
5m6d6O5b0wKGSKOIatQRS6qyr0UMuT3EbIjEJ+gg9uKHzABUAa0bZkebTGbJYEvNjVOgxgFT1dmQ
upmWNgCqAJtchF8Sz0ijWRReFdqoHv6OebyCzGeFhvOsW5BVWYMOoTWXKlqCyGe90Ov5peAqO5EI
qeB4so09WUBoGcPR9jndCvyFECQfNYU7615t73jp6gtapa2l32Dn9sVVWD2mYtoHRlKCSI+2D3k8
fDTeOxBZP3llhMqjiw/xFJErgZcxvPY6vywBRLocNaJQ+2mSAWPbAbSMpplsjnzbDHGcOAITaD4v
EihbVaje7r5vdZp+NEVI8/pPWshtRCUcyAOdnz4+0g5vgmey08qtqT4VSr47Q5rgcG2oNYlsb2Br
/mlJfARKTpYGQbdEgnofp12QuR8ZXQsvo+BvjTDO99DfluTTC7+s6tPSeLR5mSyJgaga84ULfabH
oIvN+cWa7zHxoOgj9yABcHMDUsp4UcpPrt02Vv2wA2oSR5kmMTJS8jTSzOXxmhjDvHqHNGeD8yY1
zvCHQapx8twqjrMby/7ABLhXqNm7QmdApZFjIgXpN1lOBeNv0HVJ/Fw23u4eTCqYvrm6WHr2OJ/f
2Kg5vdrzs8X28h6htQQzOyj+5XsBT4JdcAs72xB1k2TNa3Yy1QyIbgoF/MXHbd/SDgEVvCbNqA1J
9eQiEJtzfolzWszcm4cTXeuCRlOxFTT2aC7TmbFPPpcd9lDCQEnYzThTxCISOnqCTz4gH+OIsSgT
iBcYjJXboq8FtHK7kUWbVgtAyCpAQasaZ/97pLX72SqSjLNjFaxV0OYdCLgGYznECGaq2UW67rXU
cs+O3kIjMBNESt4VGpbRCP4LqDPYC40XOfQHLqCBnmUxtUtDFt7oqqPs4SYTYBDQ7gwVeZA3P6yi
9vUWUGoIbwkP3OggymoI6/11hVUJkGbFxaqKL0N+OQrkE9hzEAsHede9Nmuq8ED1Fpvz/FT7oB/H
0EQR/XXlLrolvbtmR2pmCC5UlOikVlIwIMBeZLKLySezT6pyvz36SRVl9o0FbN2l4P312j+is2QV
91qLA89qfMCEycgKLH1fOpa7/zYsgIBuZgKZ/IBFxB8kpEsQBnbpccFh72zfmpp6kNfbsxpohdVj
FyeQpGj8QPmzwmTzXeKitGvlGs/oEmOxcBIPz4Gv/v0e0zjpCLE0A8zY9y/KgBaqUHZszl1H1Gu6
TzowaIiYwo6C24MkPoLa/d5qy3lsQG2u6oYzCveC9ndyllf8Pycm9PZs64ucx5HRE9pOLdLUPniv
YOwENtOBIW1IPXEUCa0zKLzyTC9t2ssYXrztBhFt//L5NabbWzg3k2GTCxDl1xXnVwXCDCFusGOn
0Xv6vERos8IYmITQnRWSML6/fvL1POMCoYh7ebVHuTEkXFAn5hV1FZktAhSUSJkycywNjpE5YCZb
WeWmqno3Cnn9RGik7ui57urtir+5btAQWgIZCeA89IKqvvyQHsLaTj3ZMo6ODsFoSNcXgufovmNZ
fPoNf49WZhD/OoQchJ/9rkwe4Ll8ArWqiPIPAJCPPlscGTELMwBEy/R6FqQR/wMxI4DBFBiN+s2i
QkClwu+griEc0l37bR0TKN+etU7l8vJ8Xc+Hv/bLMf3+MvuEX4sNdMijq6wF+Ku23uU7JjdONOrg
HQXVi3CdfAG3dqvNcSTcqBs9Bz9ftS6ghiydNVN04/kg8aI0XSoQIqlGalCFxV8LAFavRFcJt2H5
da8QxTQepElI7Me+HmCPaTRJcULdBcSIZJzzV0BDOZxlA6mPSpf8tSAlk3VYZ78sjkKlfuB5tWdO
ZwVyjOyN9uHTt93f6WmaoR8ed1R9ugsdOrq8AHUZv49+4fYeah//hsWEWptVyLwNVrp+bsV4K6Fc
Z0CkuBVckDu8ug9iw1QGYDt9IsPKRuafo3B/KGmJ3vjQH1qJuIHErcNe3BIoC0SETkzruG3HmLDm
++w2GgOsy5KcLW8yF5J/XZaaIyMa12QFog0icle/7/dfIorh//YI/SteFqoj3LBpJke3pcEAxFTj
i+6CfVwKxQ3AroDxopgJrXr/e4yTrkuxMk99/fjuqlWmcT8PI/e3u/KELoRjhX+E3ASRyMl7Kvd3
lZBPwNzT1eJVg3VRDaHKzvigUm2H92hQMd0jesA9J3Ic6jWTKZJdenEvGSNNho4ZmRlPPAXOzr+0
7jTSvUNhqFDYWcH9ELZGn1gH8AItphtwZuVt0G2ChkUp0P9sfhguVsADUqbi0oYxnKox3rozYrIW
PibPwlgvygP5osENF6yvk2YD/4yYgAGsIa2Ykxy7Y7V8u1aAc5yvepuO8c1q0WLUMolXVzrZa4yE
A5oyyrebf+Wiw0KtH5vfft96WQCMEHTShjdE6ZSokLjAQyxMItakoDzbQDjWQ2PDWv2FTHRsba+v
aPmHMZZnLOLE29fnqz1R4HbTMIhZRBSz32ZDfJYrEhiyMlgwEi57mxh8KtGr6wMQ7uB0c6Oeqg6G
eJZ0+Bl93CfVyXkZAx9UL8L5nni9ir7eXBtyvfdtUDIc0xhHmqyvzR0LrtjLKF6rAnv8PWS4hjc8
gimhqe9JFSG1VTOkogpvbMCaWD5ded6LsS4fLbQQ8ns6+G0RoQTYbree/5Qiuw8CGaYsL/UJQroX
+VT37mzWbOTt0mILKHFyBisIkGOmO19dw5BVOUolF3xw0b1PR16LNE2uLELfc3mhxD3nlBjL5fvH
78bX2JgAIpaCzuS5XOYSiOu5JZhBn3oD1dXAraZF/UUDyMTORuEsts0g+NfUWRlMCSm6w1FLR2cZ
6lM4PoWuSuQi8LieDN82ZEmFl/3RRVs7TbLuoAvDoy+zG1jtcvdQrbB0kmCVV2ED1ZfI8KG4wTTf
9Czeexe6IPsYbucrDjCa3w/CkogEHb0vrj77jTBbsNHwGmitBVk7N9POn4UvwzsFdlwi9GBTKH8X
U+mCHsdCxFD7jtsNXIcAwtYD/+JqIfAhMw20TKJt5j2sSocn8v6MPELX9MhwyTqOejDGHbYXtc/R
Ie5MM8YyKKUl0nkPbUFck0bMgOHllGY/Tl6e+sdNSiZDFN7vYvwHWeXkNZclHAXCje7fpAxiNjTX
z5gO9RuLh927VnMCLB4cUmYIpsJUAqJHJsMhVlSCn5I7wtvYF8/GOfYZoLUQ+lsz51v70yqbTiu7
UXBXZK0osR2WCmt3WsDK6NcHDJ3nEqh1hEcnVoQ/QqS63QYLqvTzD0WzO/eBBZIYtU1TgpcBm+FL
Rm1LL2SoP2DC/cr4UaJFHS4ahnu6cevNCuohkaiOGO5rSiR8vkl2zotHiP7tAUcYR/Ezxp++x950
jcLLo60FjCIoqC3U0/OZypNpp41cEarV9lIfe2ZfRk9KPnotn6IHbGTY9HX9RumQVgNvdICaCY82
lxQABIOy38kJ6Og5qV6O/3hltNdYwbxDv1XRd3WEInXjaCjwoq3hkOKGecSsixAIQIZtpCwQxTm8
4t6l29nRORZ/NphXS1qV98zXRZiQHxBEiSqhxFAWfdK13ok7agsdst+N753b6yTyV78mIWejt2JI
UzblSBr0y592pIDJhhF7xhrkBo2dXksRSFNksm97sM0iOMhpgsnC7GjX1G9jRNdXgim5DNAElRjZ
6MFhyAH+lMhk7WHPPKbhVq+nJCq2nKo9tuhV1FbP9Zfqne0jhMpwpMl16tEWd1ejClE5yx94qzNx
33FV2b+BW0YbOXRbMfl8KVPJ117dZ7GxHfzvVlHDgO8XrF8Kymd5MoA8fO1yckutLZtjNTaDzIJl
gTId9Xfg4DEDIJ5Js0O5s3xSMI5oN5IUyyhfmsHEXaeIiHkJ9k26Uo/VQZH2TjkrNuP5DTc+WN5b
Z0Iuvib7lhewzEr4bMPrO3xUKP1nTh3RwZYPo2z/td4zsr3eLumZaBqN/1FTIhjIVhhUat/OrDTP
tOjSaiqjH1PtBYEVnbl4j7t2+BWvY+HtUCKPpkfcNvInkqkus8YxLO99haSe1HP/Tfn0tAIUClJf
zk+sYZph612ddLPvOtDKAYs0BA09D+p9khsE800jxvnaYQd5pR/b+83ohtwF2Z0PKyKrEl3bzDxg
v8gvPnQZcDVHnLoqTFPdB2GgwWDBwuJBy51rq3cGV2GBOh+5SRZMfl7U4/94t1AKi4Rfof31YQKy
0VaKxG1Xt/O4oWDg2CX0qpGCrF8IIV59PVUMZQzXenkG0+lqSKWAVIkmM6CDXFyd4VfOGhymkhrQ
jEgPaoGIZNbrxKF5YtivwNGTtBWUDJ3XaBgVZIwtJITAGTaKtp62kjvLvpqb/843KaDVqqE0Clp/
JGmvfnzUxYUe1dkpmuhT69CkNP0RtMzDC0UOGyJMKQDoCc38GBFJxO4ckngco8u3lAfLxmT7LnDN
8SapfnCLONwfBbz5izm6gPaFzYw2mR/kqc9ve8SdtG32lusstf7sNuJW1gLJvyoRATF9euw2PpGp
QXgsYHiok/fOvlJtq3SaNpeNur/apCxv7LXQIneuK3dorCgiYawXO8wPpJoseU0GJVreXOPSGmez
AAxZvo5nliIiP4npW2Dy6O3h+1jYh4D/wcvqUbg0/1cW0n8EnLha9x4hXlQ2IKMsnvaeqk4Yu/Sf
QIvbTo1qqXckO66hfyuwU8l+0mGCkShxP1nhOOKGSVoczQJsSCmOmj+1jYq52bzK66eY7iKIWlwQ
VNTzTHHeipvHs/mEVX6orfNKWBI5HcNjmwgv3qSnWIvOfHjIV0Jb8bGN/W2FvI5v+2O7H41Tkcpq
70pTzEf6K+q0ZOBQXyzsHRUcqyGvpHDph5hiB88TqIQZooJ/CbfBj7OuVOROBESAuGihXin7O3RZ
40bz7Zrk5yy2DtneCerWWX44DVvjN/uYsOGuv6if++msIT5jOCyU7bVqt/ohOpm27xSNduYNii1m
bvr0ZYnDp5uyvjZ4uVjBAYH8TAFheaIiE+CeLcQ0gFUVmWV+u9UaK3o84R7ybyYmKT4ZNbeyG3Zn
z+XgkrNufNbLVy7GTsqAbD8qRY0XdsLmlsQS7RuSgNgC4td7914HwAjcsKv/7B8A11kTqLMdQusI
nhOGdpSgDPssQzh+FlrqmqgYkQulCNi0VRczjxThyiXOjG6wZHRoD82MB+K0tXbAbOySLBcApHND
mEg3RrGQ9UqWhSNzNUqLdf9zhxTlTL3wL1Twsjv0cZqowx7qWZWutEBE69Ro8NJo5/r5ZuT2bV0k
sRS6n14JQSrM/0+8uOGo6zZHlkar4B0OJ3Iv0SqaGI514YUkDxPwFxh03+z+N7YYqeW/Mv23A0Ba
Wqgqz7o0nbFp/R8VwmgcAga5YjVj3WulBlEL9p3lbXWNNsNf/JuivzReS4j/kHpwgkpvazdDkC0l
miCUNWVGQPGFBCVRnnvc7KLGiYFAwmHfFAnS1mmWqP9lxTNiYFZ9hiNv6Adf5eDHPpUyLT8DPjME
t7CAS7iVTkw8q9Zp7o5ktpUspqcBmtuR3GTlR1DMAbvWv4TooONoKF/V0IovjQ10RFaV6TWotE4n
caWQzWbe2tpvg3WvLCz1Pj/0EDcP4gTcqPG/k2ItP93NaSo3Ueb46GhuQXAFUvLlNs3VDnn5OKbh
Daa36KrC0loAnwhBwntcxOY4P2Ng/EyGKOVnaGMOktMBZobOEe1ktW8YzprLyVt1mE8oe4vWFHnH
dYKBtIz01sZynj5lIlJPqSfXVDTUTioVAmhHAsx7UJrniBoL1QqTeEqOfr2Arir1mK4N00HULIt4
dyTDeEbZhTuMN++juyLM4aYY0kKBsOTEKSDnUXl+izQjth8YCezF1DsNvtwEmuW8eRqg6VIU5UFj
PxsxS/5QyYa4LUilK+RvGtdp2AuaxFKUWra5nhNp3kGzS7y4cTUzKhNiZWoDVcFSYLPrKq4fDkMf
PNihh8QdoGgF0TjB0qxVtrQFK6h0KlTH/mVaG1lrNBM4wzySTwLwhBbDnZMaOySFbe0DCTf20tcM
siYQJptjsR+EhWhQzaCbkSre45UJ12bVW7Eo5bXGwE5KHdYlaPaM9DcotrX2cHGxOWGHfxIGU1u1
QEyzY+t9Xet/lWlE1tfYMC8Lu0t+zRXCJqNsMCxel+VkBuuS7a02rbnFHLB3Os/D31LU1U+g48jm
ZMMHfMvxT5KtsPNbboa1SbExoeZj6Vnu8P18QOSO7DLi1o8tjB2Nxd5InUN934F/iiXex3ipMoDW
FsW9Em9QSMJl7hAFykL68FuMqqf/RNMoFgRI6ZRwMQzrCGcPOE/PiLy4mLyLsUWB4LV8ifsaBqCo
8fEGqilyVsiyjjiLbv03zu0BtTLA879yYkF7N1flkL++pl7WuOxYPELxMu0DnxpkklCDOhJ7Spsx
SZelgOcfbPdUFVEY7ztSbw6hUt141/gNn4yujD2SOLKK4OIJ5P1Zq2sIys00SYuaz6bFqxzmuCLz
Kn22CGdO1BodiOhSbhuaqysf0nCVFwPdghAdCYkMvhs/0uZ1BORfm6M789qQXAfxGgTwDgzKP2VW
VAsBI3tRDfkRYslB0f+AqToKz7kPEtmI3QW1drveMI/v3TlMozamohN+Y9qjhBkiMnLid75svujS
vYOLlEHdu90f1m+CyI0Mjmob/z6ehZ29BwapOJoZPKD4y70CaQaexeqLCTAT3D8LdsEqHttI9ElT
r3urM5KEa1mgy0o8hda6GEYrAY/NrVwYyfwJEvrTfKCp/6FWGbnaOR00a5BkiyCPfwgfRbdPsiGI
tQz+QPyI6qfz1rhhmakB7zkGcawDND3r0+awnyWO7cNmc3XXgQik495iGNJCaUZamOe7fA3piSWI
wDK2CJfcupAok25ME9UUCEOI1GbtTftsLkqOlclA8SL5rX3IvLnk/WwzimGA/GBHIMP/gamAXGQX
QPTiw1Gknhx2PEnGqNPmZPo5W9JF75ber0KytM6ZOLN5cIejokT3WeLFgh8m0jGluNtHFFvFjfCJ
t9wV+36wpiJghs9SIGOwLnPPt5SUBGUXimad911fbYVQSZXPiMt5F+9pjmhrhGGgtqILwCfEDMJP
rrwb0f6FPQe7XfXHGegp7+sBgyPketdWRsHxUtUlNnZ7ujzbiO8MKCffa+I/SxqGtnGF6G/F6UNv
0kLLl9+pQIaeoxCKmrDrow1R6+9GW+1DEWY5zBAsX+nLu9srN0h6By5nbPOG+bePobOAWTrVlGkU
eRVHoXoeZoVzxpqKNJzucqKH7JgYhsRDKGUdPh+eKA41sv9PXEklHtUo5ccy2kYo/Yfz7HrCCuZt
aUSYz1noyp/DojDIJkFyHiKPnGPOoLJzXFCv8N8mbW08y6FCjnIhTlebeLeLwClYIziFuEwRX7zO
v1eBMAUuxzUfQc/v2i/MfH2JgIb/vwZaXP3Bkc/SLC9BdKMCR6dkZEtc/3a58D5RUhdfC8dRY32M
XBnqBnJyYSPpUPu2WyZr5lcHn0XAdsF6bgnDJwxrpJOdDZJ3zmnqbtbCo4SWA7yIEXTRFaxE4HKg
cq9D759wK+nCgpFR2vi0ZNQ5s2x/v9Uubnu3gIbOkR0Q8dN8E4vyO+tCdWFUZbanU9o3T2e0cAKB
zt96VI3PLxnqXn01hrD+ApnikG/p808pfdVHc1OEOKboI1HthDLicpSXvH+ba0fZrocZnuOD6+8X
+P/UD+VC882uAYv2kgorKTiq+luy/x4/E8SVS9V+wA0fLKuW4SXZP0VEZu2D7zh/5j5haeOYzOIz
tcuEHHDZtP68ah/unmaWZTMjSkgOZyCcABUiZT5fEKJ8FNPt9B3r2czm+Br/jCfd96XWr804jyb6
7y8hYyygNWdcfkTFp7Kt8Om9iAoZVXoQItxNHhS341eTegTa9EdxKmqBFIk2EWzKI3zdsszwwDII
XbNnKALrsh5V6Y7lVgr+iLUVQfF5mGxAerUQgrGDuY4ytCRinozmWgnN7tiRGTTXgUm/ilG2zjAE
2aCvYSznf+1v8miwwXbsO7ggd5qVWveP1LBV8+bshL5LVP7ixCXb8HTYTkOjhCUr9iBipQGiCoBb
jt1a8nX+Y0WD74S4D/KdK63oIb2gQZq5JXi90ovoSCHeybZp/K8GbOlHyAmpXyAP/KLcLAa6jpj7
cD0zvjVpNAmaIpj9avdIGi4NhBGKQt6pmwdaVQw+Wb+HCMyfOCMkiS1f57v9ZEbgpQgecZY1gCeD
vaDj3vbAX9sZuuY0zfxzLRw9mnnDTE3+b1VNRXPDE3Dl7lowXQLjfY0+r7Y+gir/P2yVeHYoz58s
aRPJgD4QjafzXVFOWIJA/oxllW7WhPybeR/tF1pDyu/YxZXelKmdnmWUJLCbAaTUVq8zH5sFGVc6
RMM8lG/hgE+84hVL/XiG+xgDb4wkTPX1RusiBH1KwIam4idbhIrOlRn8YDeQ01PlXIvTLrPmST/Q
VBnsoLKK5Cnuz9CiWc4bs4qz6mKfT9WvStDSMuJv3W5AKEdsEVs/P2+f8LHctN29EXQwSFDDmkVf
QfKgwHk40UyGazM/5z1KWe7M/Ofus4exzCo+hdaX3J70ra1pAZhXi4tqrOpamDBq0qu5fa5/hXnC
yxykT9tpZgN3g5SKf5RPRrTLwoTdjOl1LP1LSXi+vKz3fYoZvbuhGqJr/A6QujQC6/pzAwBn6r2r
sxf4KxnpfL4L5kgGXtveonEnYH2ETTfIN64YwkZ2eJoTcIxah5Dl2Pf2PEGX6zY/3XEkhbdDxSa5
G8fHFc7VH4kMjs8Q0ztehSuFkxOtCMYkytcgPn4cuO0pvEhz4HLvmMnTKio0MPNJvv64BWoTbduX
ba+689HbxoUD4ADJl+BCw3TdksSxBnap68b2vag1QEkHm7MmXr35yMqmPJYkzzRWfBP2nWSgYFWa
7lnyUQFmx+Wmz1C/G9w3/Lx2De1ZNVoO0lktFeSTM+8lsHderjjcueIzQCa4HYDADsYvykc2pWjq
R2QZ3dmE3oFdDhwJieTRgXomoWY6z85+6mCMfgHH5V7u+aWYoeQRNt+HzancLy6i/fAcoMOXBp5S
+yWfMXFL48kbDX8MiNmc4EExQIcAfXBcpVqL9clQ7EEZvstCbquwCG8t32fGSzSnu4GV8CdP9ITB
WGhlvlCw+VXwBqaTfembnuYFK1Impi79L3Z/YS62gXkazmFhh+Gi/n98qRiBhqLp0DUGR+sJ5pQo
j15aa3Bl8DY/Ot2jnnRiIrLhO3APxChSxufwB9TJVO+bVKCnH3PbdtqgTmwqu4NBOWYK7UHsmcKg
J0+g5J7RP4B2fhG8r6p4T+Km/0UuBJWleUXBz9IiFj8/HOkyxrh30IJ1XiiVlXMjLuP/51x2SiLC
uOTZJX8xVcc08+qcxzVWp8ywvGuyWTsHWRbrUKqCDUJvNBqLqRzsSEr/leEKh43K2b1y1WhCgvTP
IUyYDnRPZX5ZKAmC8+8J8e7p0DHkONfq9AtqVyS7l99Gr2tzU/2JrRPrzNeI2vECLuKXam3/HGCz
Cv03KeCMzkBwqHuUgyKwSINefBKAqaJEDGswfi8Dz01EEXFsfSvvdWZW26fYDGtms17OCBVxsdt4
YCwu6GBl4s4bOj2xMD4BZ/XFED+vI5AAdT42VkpQvHLYtvaGRGgZ5qhp+GHKxQd9ByEtaty7pcq+
+QloAmznsLXTi5ebl6Mf1KT/wVoyuCfYuacRiHJ8BBQSqnpUSljPDaw1K1vDzYdoYF6Bp5invA3r
ZIGXGSvmnMCikCIIQX4mNIYd8lcDgYBE8WcLuKMROpKQOugVwlT6nGBOMXKGAXbGKwBMKomn9wIe
1EnGa0yGpD2pkDoC5Cl+URxhBDlMiGXI+iXow3sxcqQuYGkQBObQ8Hjq0ej7N1yplEAlDXza4REF
c5xbiqfE5fiK5Rk0TpXopCRXVR4/R9/LlXpA3txA5782tmXKX2cwaAqoAsokc0/H7LFe/zZ/4mIM
Jmdvcdu3xt8OBQSu4IOSZzPeesuCThHCRxwmi4L+m2tL2gPFdBZvPNeeTQbLTMxm7g3d8gXloVKT
q+ptj3S9tfXwzR7YjiqAP0ao7oMTwAQeJO2LDBXfRdNXQQ7rLunBIwCy3rbE4FqHNPI7eQP15Nfq
8dckdk2EtTIe5AW0T6WR1S4kRHglNhTp+UATirasTLcUN1fqdap+fmYHM1hx8OyejoB7NNjBevoB
gB47GIq8lVlpJyoYn5S9P+xaXVvTRxCrGl0QK8/X7zhHEOWr0r6mILHUcTiIliGhLI6ypKGCKcbz
KTeUqzzRbz3UbX4f0yhcCQTB/3RYjOcesbnrx9kT7zNnek68IJct0b3k4v9W0DLsYCaiK5K3ELHV
ZJK1A46g8mIXmiAITBgFLSo7cd1gOgI4IWusKXt2pMe6XjRVRh9zcC9G46xrauhSMKbAIRCNF9OK
U0b9Lci0oiU16rqHxjVrBlpi6XLZGATUi+DeCWYbxSayG6IPTWaIMwmfGboGBuLUcT9xgrO7zMFE
mt9LeyBIZphf1p7otYbIGsv7Xm59Nxf2f5nf+pBPltJ8gFEkW1PKF3hqCY5cECQmq6gQOeZe3ZpC
UpbqHt/wQFCmwAmXYZq3AfmUqEUiE7VkYU3DEkntE93qfsdre2kLBw0Lg47jFUPgmgUdmCA4hGYw
TtHwyQj24rvcffXV5iXjGw0nMnAymcR4xo3FKgAeSR0bZIESqnugnus/OUSRxVzFocNSFTMZg8yx
D1qjO+xZjXSTZInQkqSj5bHr+BqbsghAPxw9PCw9qk93CyE86wp0Xwp+HW13urvOHrQol2jEZIpQ
Q9Sloa3cegeU2Js99eRdK/KnJOXUryLfyl85UgLV+zqV7e3cyJYObnk9QzGXCj5B6eNq2z+/RtMP
GwB8XmKzqqGOdmblN7juQmFE7hbYeV5JTMFxBp8Aac5P8uk7iEq3wKwJj9c+NmSRp7C8pr8M2/NY
3nJXSSokarW3CHNWvouLvD6QLfnANubWQvvAmEKceUj+Teo2p4+OYdwRph48RPyHXo8kaDJrBjF/
Cm5Balw29osEUFObd5KxsA9a8lLAfw5H53FS8InEEtfPJB0YcXOjcgOoiOSZdAS4nqhnlc67G1fc
SCgfHJs5vVT34roYFQl8fmWTw2WEuPIxiMo8PWptsYGUD4vUBLkxQ/hT2mhSEkzGP0hpAFjqe6RK
QJrkJm+FbS+Na4oOjVPuXfq3ecdGnkWhZIm/GpjEu6KX8iEsB2y/X7+14VQwk+W64bvaCvyIYfw0
pCICItGrIX3E2fZokAWbgdVSV4d+a60MpXcTTO3Q0I8AOp7CJq9IO481OiRf2e4UaUmZdPrsQzCC
EL7IVJS37ujEcgzcjyGnzc3BoQlmIcdQ9UNns7TzttfHFP8KYn8OYlIogVmhbfgSUfLmrzKlRAMk
lxxcUcpKjMlsj3o44IMx5HQDZeHK0Grv9tDXBgfe8fPDrrvu0yfNpoJTgyVxZjWJK6YpRHutQnr5
j7dMNxyDRZlkqVytXS4QdGB2HlUXqPJlRMu/7LZbAWy2CaS8Aw+GbhTYlOG+sQh1kPPh2geNPUWe
Ms6ir8JkGAdfleTrVcjop4EX8DthO8/zATdpi8ViWcv5EZTEvkKr8CjNH2R3MyBIpv1ml8KKc3eI
gN4EYqg537lIKEM38nc5FcQz4/9dAccaR2bvll9ZOOa50Q84Znl0UWFZukGULVDXnFhaYng4gt3u
eek0K9Xy4x7KhjUOpA0Wt/maQgQl8Xqzd8Dn0RhLxpy1HYpSGB7w+EdScJ5FzJYKgLnBDZvkpXZ3
25Bh6gCzYmfNBlPLsPOpfCFh99BCcjDRoF3vv2vcrwdRVCgny1CKVR6fgIDX96DAcMWnLr+M1/y3
sbLLHAGz0kyxrmjxtLrfyqHE2pvw3uBBC+4l/xX3sLZLrVTAL15AMqsXzu+DztvjI1nob4vh2hu4
KHABxcCXXRP/Wn81kceo3U2f6xOaNXEoTKxHveQZV/iXii+aVo7U2T3uqnoPHnOjIRiEGG2ndwS+
FJhdVTunLSeXN4FI5bPTZb2REGjrgfDl9qPrID0/AcF69yS4XSYwgfKVbPh0F0cWSFBqOhy+WsvM
k1G7hlzBkYWf0iURquKD+/WoykVpebCu+j5Qx7VR3Iwt0vS3pLyfPTTvMwE/ePuBGaZMnuGv59ml
FRSffwsSTr8Djn3TVNFsi3yNoyFPvz4kTOc+SOzfWppmLJgnI73y07gbYBtwtnYrf/ulsly2kfVb
aQMZh3Nrdp/RqLB28OvjPqFg1+aKtc34EaK/GIFsm9wt6JVx9BM/ivwL1kqj3rSlvakRBWsTEOrI
nW1tzSBVYlr3ozWQ1ZX/Wu4WFjBuwtcfWE9n8c7J94BOf7kVmUHzg8L8ThUU/q9UneyjJgwTuXnO
z3P5u1y7TMNazsYp9HQ7h2W4LL1DEfwqlZBTQDFR1wntXYoHO0dkPqh+cqrUqCF9Tr0GJbv1nVHe
p469rF6IXK7v96izYksJfctKXR7sj+zVCDl/s5F+xUKv9B+aBvnIu51n4DaRGZScky5YODT8oBeN
YIghkKfzJ/88SzFenVYPlyIeIESg5pT4334vf4eIGgXZ/JN5noddCNuveYmCbqdXDPt1ftf2EmrG
zimCDVxBUOIAIMXg/4Uu/HoMHwjqxXh3388NpH9YdDcg58vwMoPVYjLPaMKTh/XwdpTZNQ0EYlOg
9lf+7yynlU2U4WrrGU4oBaHMMVD/zXPl+ESfG4YJqja7kmo5xNde4wdXF5uJfgUpr+ZQfLh2rnnt
FbaGpkndnEq6gvO3zrnhY/wxMlT+QrlZXTvSwy3Vj+jVdzOvH8I+9tkeJbqIz5VZqaACTXr979Tx
zZy9s0vo+1yyJ/U4fGADvTtULiErtX7+/igkPv5Ts9qhUSk/RYsTFzZgfbPN0qJRzOqn6TjXCk4l
4F/eSj7sDNe91IQc0vwOIXlAfGNW1XGxo3j3UCvG+IEZvfOfzswxFK0mDy16CS07seZw7niBPn3o
MCuEvwhIQPwUmEQFo44TmnPGf151VvyFqrg+KVVneXZjtw/2cC5liiKmCpDtF1xl7vs7vKlAxO6J
VkNOb8su/eLuiyLpH91hz/Rl8hItU2kMx2G33Qh2E0ETpFzJtnkA2ISPUqPqFg+9N+d4qzplQ8uU
nqwgPFnTJgRH2uWA1gpemPiZmxeG3WlYhw38wZSH+cJPYmC7/y2bxsFy4D4yqqtMgpkIYw5FKIWq
w7MMVa2Sb21W5UMslMGB/qM6ZJA++PPZDhhyER9cG38AGNlRDidUCQzkwo2A0HA0FT2ut+QekRwh
kH8WbD3L28NJhIuWZBQc8CDDcqH1iToshbR9jObQF3N92OBWCSzZIzOIv6qKe6N8p22uuykiCMIn
hUd/hTIq4AY7rp8uaqLpQ3LENNVKglSRaNRo7TcJfbqiQN45eIePzuDtuLp3yvbzbbAI0ZamO4dw
5dTNOkX0LroOHH6/SZAsWKhfQjH9k/QnBq6Zkhw6jgYQzPpwLviWhKXIe3F3d/M3ov4YpZTkU37h
Qan89xJnBT4hlMk2n2PKrYBCoMaxxMdPj8kVGd+gEB60gPn+3bRZUszTOmVfGhSIeHK93paC7PaK
rdY5P74AZ63aWGr29jHfL6aPN1MOjnte8oe1cAMfHzcj4me+XYIcK2h2hg0qPRz4X8VCP69zWqAg
FEC9yeeD/Q5b9bRnEvmspZNHjqEY7jm/oWhOe8jMJscp5t0YniJrs4wc3J7+4p1bkjoj/o3azipW
qiC23fQF0/FWXrtnGCMlIeveBpZh8v/zl8OtYQ3fSEawF91s1GgbTSPRVpmd1Pk+B0rhpOsmO8t6
KYWzmB074LAbGjk1O6JhUBspYxSArSwsvaYmiCYOParrjMcuOVw2D/Lc8XDgfhRmHExVf4bH5kVB
zuWLlk1B7vXmTZ9XOEK4YzSGneaP6BAqehatTUyRTWW88Rduuw5oW8syt4Hw1dbx0IfGMaJzhnY0
28GAZD/TjTqSC3R3JQ0WSHEdnvHsYAkf8MOD7JuqUkqN3m552Wp/3wHwv20k7dsfvV6xpHU9S4Ll
WHGjqo3IHK4WYeTEDx5VGac3Pi9IAZeptuvcKnzYA5mjOrCCSyQT3Xpnmsd2HjsudkDMmegMF3q+
z3ZIdXCNm/gdJPB4oiFhXGD6oLfBpp/k5lVwoQLdKX5zsu9ASgBSEOEx+Kf7JW5nrBiXH1YJvkw2
4CZ9axOaV8tuNk7hNqcxg6DHAWHpKYTuvd6GMj5l0nQJ2YnBxl6lAkeoo34ITJnyYkFxpgu+29HX
5sMT5vfvp0j+tUs86l7hLyjs/KEwNzSte47yeYcflUQeywRLQ9J1YV3BENfBlu4hSxwxEJ38ehMN
jYX6nHBv0rUpGwVGCMWzJopFAUKqZjtn08oyMzfYvjMuntC1M/m8pH2170h4AoClZjPxp9qklTk+
NaVL0uuUZW7FsTu/kzYNX3lqW1Xm7qCU/5pTWC2vqavRr9B8xilj9YTVx98QtHmSRYRFdm56YsQm
xuRxumaSIp536Zak4QtCVj5a1VVpww/MdWo+xYsKf4xjhNO7r696MwFeX5RvX+dYhHJG7+FRFo0g
kNShlMCqg5dc6Hr/Pk6Xtvt57Q6BJ8xhfyzvSkLTPlJwd5CUkOSCFcPEik8flkKV9Yg//dNeCEE5
2PiZd68SsCeBvQ6WveA13JRQYMWZq5ocVQqQST/b5C3x/jvgineDa0HvL1gTNFVX6X6uz6DzRN//
jCvC0v/oVGoEwrnn4F8YPOTEuz0MLCtkJ3RwEoFm+9WH20Sw8NjeXSbh/otAUjn5rdf9vGDt+vtV
0JZA2exOxQH6BZc2elO/YUzpAKWymHwG1kdIdhA/P7JvBtSxu/7jM6rfy5s8TFbDmdHS7jMWsvOy
BBhf/bW42cNLFIe5G9LluAI5sNdsxspkWeNx4FBa6R5/Z7vZ6A0swowFoyiVXS1LncegymYz1Uad
B6N2Cg5sAtvuUFQQHBtRBSyEt5dR+UWX8Zzug3gMIJ6b4RUfLQskqt9cLlnRzmDsHGhkh7+COeBm
wfacP19Fl44Gl9ugXTCT6YdzqXIP344swcHkBQkR6raveAyVsD1R35gu2OrKwPOKXvGNqDoh2XrC
r0eXMJxODkpo6vOVqQo0kUCkIoTVEuH3y1j6GHFn06HBxWfloH+H8w1V0ccx/1qoersBAMKSK+Um
PmPwdhWAJJhLTHccI/S0ceRosC5VtuNQpiEtQbZLbX8FQ0qvAyUf+SosZOaWZdtGWhj5bOHemVjj
Z9do3fylJ2K84X/TD9WhNs81s4rhERykZI6rEC9HLc7KbStzRJc/vlPpaod8E7NK90R6pA0pHoI4
kZCrdNX/bmE0W0yituFhT1IsRrXzS0WcBh5YJHgvMprgPEhpJCvcH546WH/DD5PjAZnSGw1kUUMg
LInCMd5EkFiRrGkqcwSE3KQD5vkIKHExBrK/bo6jfvNHc1SCHTX7XM46iSNhYQbExeMthumr+PoU
ZXgf8DnOCBwy7bB5u4tQATaRva7EzrWn8HIHwR6bvSN+8GCtaiwsUSODMWgsck8Gnod5ejhtWu5p
el6bOh1hM4JUvlvKdDqALHjMnGjNk7pLFn4Jid1ohoGqxAjN2ASJ8gzuGWEkV8KlEDWwRK2WS85F
eCLR3Pu6huT77O1FR4G+k0i9drJBXewYcgdndyo+SRTTBzQ0CXlHuHAP12J1g4YDXZeAoxyuBGmu
o9LPW8cDHHkWkRVLJrgMsN72mXhw/Pv/fFLChRHWXJs+NNAQAIEEje1QzhFG/+Ossouf2Z2oDlb1
7GUq3jJy4Ftazu6uPoqiA6myhAxO0I1m1apjDf9Dlkrc0YZ1sDQY8A+Ju1ZTl413Sm89y3zO1h9N
7Yjraum/QDkLNrkwsczHvE7GxLSJP6K01sp9wNdT61Ioi4zcnXMhqezXFicB/Cfso+9p2aC/XNzV
C2QrS5f1LbI/e9fN7/tIOz//UJZ+P/v1HuLdF8s+o6zqoZm4WPbvQW8suhKiUk+D/AESmE+HTu61
DUCPNWdfpwBYgYZ4xthCWMtlN7iurJgnAiwnTeWN7pY68SjevT2hWfe0+i0YFuyOMaZAvQL8UChN
C74/WmzrW6l1sJX2Ukdn7SjfpZBhAWpdJW8A1t6SpN/nbIyq4qQOcb9sxGK6l+R/9xuoboioDuKa
H6xh5bwavJu8ca5PnrG+cCYevvdDH7witBGV3kOXqQjnS64fVPKO+9B8HZmymtu1T5NojW2+mYli
cjyyc+nJqa0d642BCApMzxhfZ9peVN92d1RVf6vH63raJvTctlgk0/qPLGXxYQEMGw6yhP2gmCfr
JtOvdM43KgqW6yzk2X3I4NEp6hGHXEDo0MEy5UB59SBsiiCv7KZ0YnKFhVlPoh7GCOCpjba/wn5b
SrXcxusAMmc7yblz0OdlksD91lYCsFz9MUSsbN0H4+T1M4hqtYil8u92qCu09A7QWqeVrFS9QM2V
+YmRf7NW8v+DHb4pWTGR72VWp3eU4xKFga/xmAChYDtc7l+S2odi3Zad5R4tle275FwvBmQqfODX
BatVSxxOZnNOhRLHhRte3wza7dxBb+SQKdeEDxMdXW5ofr5+hL7DPaAwEZSQ33wmXaFeUfpB8rHS
QJt/qvDsnrujZ5njbAo9Hm7HMUUIdSjsohWl6fCARKCPV+/jLAt905Bsr2gPL/ql5fnAUjC0KEA3
4XLBDiOksGoPzHO7Sfg1MEq6k6mQ3eYqI98x7EbBSJsCuKJSeVeYLCa1vEYMhbWAGc7Y0pxCyw5y
x7IAnPpCif3+gUZiGYLr06kPJak5rv9Jyz/2wvAJHCx8BPKih1gzFgHmfxIV0plogQjYHoEUoyTe
2pVM0Ss7ZsnJuOUQPonbh15C4OXIWlk9ZcYzB8BqvLJZDKGXcjHJPfccJBPpu4A2WASnKDaNzzAR
B1chPcfKp/wQvdmMjgIPBAgEIlHIWGPOBxuSjq0TYMGDYf2pe9v7DeaJF22XPpxXh4B2tQ9JeKFS
BLrU+V2qM9m7Hm5430aqNdFtQVOQW+CEeLlSy9uONwVShEo6ZWgn7egyt5ftNPb5EMmkfSiOGenJ
i7QP2A3Bwlqhk8F7rnEwNXNVBDzbFWXLevk1TJ0y9cRdln0EG3DJ1FPOK2eOoEvN1Cd1mP1F6Twm
pF3QFdm4B04ruxF1hLx/nv942Md2TKYKRt0pk8eiEcA7U/2om6IfjXFavyI+eeIPxnvudDvgyltY
qx4n619VTDnSTsLewuJJRILOWm1PQhw+J636ehAJowd/ni42JUZq+aWMi0R1IxjXGTk9zuXhF6kM
XMXwSjIffj4y9LIYZetS9qi3SYTKb47V4bC/tGDqTNkuWxTxbRlLWIDn308C+wBAzYxgaZ8XMNGq
qZIrff9CDrt/+dJJ4NyloW0/N0QDW1VLwvYofmP1bioty0wjbm9iQLA9oJwXRrQ9dmtHVX7aB33k
yBSeeSYdS+1uk0u2RHIkN8+DLrK48EmlW6+85LpRyEVUyjpa2kF7zkzIiUol6agGOTndPCVEhNhH
ExUX/gYfKzw6ul4DS7mUuE9JZldpnP9EQAxbJWBs82hzYGOcg80kR9i1lggi8bHYSI7JGtYgN+P4
BDUYlJJiy/j0nH3sh31i2lp33SrFtw5hYVrzutJRA3OH5B8+eyod29I+BuqdCA/Joe2qtEqO/031
OAbrqQVfyrXirqlHS9iuQwdbfg+djnFP9IsY82J42sYFSiG4NOeaUDbHMr/5Un7CbwIf35Doycbf
Btp0Eg12Phu4xFw28n7mdN215ffZ/8X2JnaNeIWN5rDvf3J3oqN2/Fu9XijEICanFLZa18qcZ9DW
ZnpeEVA0h4CY1r062s9DqSePXn/sr9iHQcahwIU9K9bCl82Z0C38ZYSiTWi+H1QHq+wCQVl2dCv4
cJHQuFeCWRXP6pmH4zj5FaXZ9Im5wYTc6f/VdMMCGt2pQyZkBcRKH52kSr4v7yrocz4X4uf7MFEY
hy6I4O/hrrJRxbKCI4PTsnG/jiMtlNiz+BXh1XmYa4K5yeLm6kIVC0axJ8LDlz8I9j4A7Q3aS1oB
mfW1YY95Itm0p61uC5sIaKVWGl6FOsRyPCJbdOgdLd7t8WZ2FcvBCN1LfnbgZB92m847AxxDIlG4
cz9FzGHta6KPF24YY2awALT1EyBXtpBhqPAQJsnAP/ucakwvq3l2jlnCSofHS4Tz6XkpY574u38+
cCkKFyO6m1gtrKFYQFlg3cjCN32jg3pZaaKpPetyuNvchj5ancX8dCdSwrpx0a9ZH5WrbK4z3Nhv
b8BIciJTXH2jQe74BKUWI/RggDwMLFazTfgWaGya43KeII19MotREE6bm43vfIBe5Yp5pXxOJfgO
Km+Wrl4KgtspJ6ey1Jl9y9ZBM5fDbAUZPpSLNUY+RwprrGDW4oDY+lBITzkODPsS3WhtX6DejudE
uIWUi8tTEP8oI64co/e7Wkpk2/42M7silU7seaLzTXFLoMy0XhNfpFK0oOiMA5Z0u8BPRK/Ld+Tf
n3qZqBXMDmgsOKPWHBaDvfPhOt7/IEVRevm+BSQ2KGdi0SNnDoOgv68VAVAbIQuzdB+oLeBUN9uQ
2NWV8fjNM4ge5nQ388YcwFSZm0r8evyUpGjzWNbOrJuHIgYPz/bThptYozasPcHGLUMKMV2+jR4k
fzbaD8Bi7WQ9j1oiumnzVgZqesBL7VyLR7k7DHa6M+Mi0ucCm8mDBAL86e730e9jRtOa9pESFnVK
uiYwiFvmdYMUpXdlarscaa2JCfUC8hS4isT3kuRNFZYwtoybyW1YFrSW7XW/mslq+GhD6q8b7e9N
pwxjYwtHGtPHf1ipuZ7HPC/ZCJl7MIx2QRJC1JTtt4RJsbv4FezpwOy/4DHabL8IBWS3Mxx6E1E+
bj/I7ki/NKO/nj2bMTosvstX1/t6o1C5Pmv4O2o7D5lINEfZ7DkbJOziyM2v0k6T5h0JzruAUwQV
rd0BrX3V7IpjQQhxPiaDN/LMGGq+BDGHf4tGVJzzMg74i0+pYiNFvrxVf9/3391Zz9PDFohdMgw6
RYhBChz6uuscDowxLNjU7taXyArjU3Gj5w0YO5n6GzhUkCoORwFHutRid8aSJz8amu719E1K5onj
6OMOKyFDtAr5BuwqzjVtrf6quYrlwu+FwrGLiRy23GCIuCOQqg5WTwS7+ucwKY6599q1qEYeHlA3
PQke3kToNKtVwvjQjt1fVUG8hF6/gguB9Gl8z4JfyNxrZnny/FlOkWOZUcJiMRq6+WLWoiXcH7ED
CxoMG5qFwgE4XQ7S4W3ZIDtAJ/dN6W4p7K97typjk2V9nXPC8BOT+913dsNihjjoAmVdB+8qC2+5
ivsWDT7d729Tq814SNjWnqr0EnmVYMaUlkdBTbAkYGURJxraJKGlIVUTpVpRbonH6cYKuxVkR+ga
q5qFH8N4c41JP5NMBfkPwnbS6RGk1IPWFHSd3qfCohWRVD6UCKDUViNAbRLOcXcaOkeQCet5Sb7+
n32G6bLNxH+y92Pn8NQuiGkIXfHoGMNY7IPpODztaYebEkJayB2uLYhHVquT7TthZV/9Sk0pIoSr
eD7D/lUGXAFEo4YAHO5DXloccdfhxBamIYmFFEZ2LYjZW3SqIuwhPwfD8Ekfk6MZUokkaWaGVTuz
AKyiiH0gkZXV4xb4+uRBVLXjH1OTXla2r7VjAVlBsk6cvOH8NrxVt8C82kCctskvBhiPCWabF8zU
IQeNZ7Lxh0iSTwhGR93mYSroI5GjlFggS0BXBgTVzl+WsqI7Tvg+0iEqKYCRdNXzra4oNjHmtZjP
BEZ4aOGvpoqcOaIQ1DBg/BljZhq5VZlObLUyt7O7IYK9iqrP1P3B2U5TE5X1k7t49QXIiQJrlIlE
EcP1Cs29rCj2tzdsrJfzPyGtuUAVsK0uoE65cmFo5goQr8vKDddFZacJ7y7ElqntFtrw6ZfRkwNF
TvEWN74hDdmKvitMwDZBCo0yN0EckVnRiSk9zW9PJuG//L/21eh9RuZilqbv4FF6YSC5iPgPLy3i
mJUwVm69SB0SH1HmQDKOD0mesF9A278oS8q1IWxg4TRNJnGKKrEi664LVftD+aGwhPFMCtEb42T/
3jkYgJlwZsIlnTUUFjhSnCMBbkcmOrtkYgksY+IKLTnqm9bOFXMou1jrNDcbyKL8lI5BOaEiLEfH
H39Tgran0JoNVOyF2njkJ3X7QDxh4t9CDyTY+SizCX5UyyneADTjT4CXEwioW1kRKJkTxWl272v6
JGhsjxDcHHO3CtOSwdosiqqujNI5xI4DdT6ghOpK4GFYMjHn+N1WY08gyMtZzixupHLivmEMrq4f
2M0Aa6uRU/oQIx+0fEWa1YTYTIgdK9fnMWnAHYMgo0XQQAnQJ8ixvPHjr8iwoVwRmQUDCL04x7CU
QAALgSZTe4G6h9njUQYF8xZKhCKBROeBt97N1FMCARRLpOlgJNfcKDXNmACczPOHiANRG/awhF0A
DKWxMhLkN4n6d40x0tujI+x+0NGe+o5X6AJUO3otyKtCQhF9tnhK3Vy4zX1HwTVoFqnvT0tJp8u3
RrT03tofQkjjrdVdKimfy37AgBrxIaCjKANRbTeupP0aU0woQHXepp+E0sPS+K/oVCAiUVlXWSk4
Mz05Hq77WGBrOPIbJOgnHmhO3iAYY9Y2sEXTRShsiQsyPLHHMeUNLhcLSpYZJTs/BmMRJcOlj/wm
arECEmmtJKCbaRVTfCaiCxm/eexnbaX9xMrxPnJU8TV4rSLu5P7BpP5HNGUoA3anBHjW24xODpDY
8lJKGa6A3r3qZDh6aCkWECLp+SKtwAXJ9S51OQwdzxG+dij288C/I5RBlzVOncN/9k6KEp5/f2b1
d/EPpaJc+CoTDIbdMrLI6LW1LJXSiwEtwA0kwQ7QjbVcQJdzySX/06xg/dBx8wwD8H7O00nxStdS
F6mCPh8+zWq1Ck7UGdbZEvnUozODmf38NsFltlTHLx8S311flSSdr5yf1dDwC0Sq37KPCj4o1HZq
BDekP+D4o4YW799Hfphsv73xRT13yA9fHgdaXc0wSnZEA5HRy9Ux+1vWBecqg/gKBy0d4LAau1FB
UK67sp8h0UGsQlj7DJD4XbeSC5DnVpoz3Ro27I83/O0kwysAlczzMqth4O3DDf8EKmX/mhLs7XK4
FqaEKLFMrXZc62N0KPXHRTIjq6bWt/lbJ9OISVL/qwDfjb2lFRqNufon+aBFD6DLiqXPQAfHicME
FBUaa2BMnJ/bhRRtn6zylj27eQwFz+69GMIMtO62ILMq3zMpT9S6d9e8dgPwCKQd1FxeFQa2v6g0
i/QfNo5QeWPEhl+dJskl6J93X/+KSoMyMwTIKcLOeCAm4lRxrtzqC0ZVpg8h2o4lZGQ5UCxPzSJ/
lxRa92uAm2lD8JXPF1K7QyDf8B9uu3vipWy39V/jNZSK9Rsfcieoh8FrFgRYrCfklvW7CmKZRk1b
sxpRBk0ThCRYVPPtv6dr1eXqT5HBIDvyqXgztNTazk2VJtQWzq74URVkJVdqfzHFfO/ryRu0ayPa
O3MGpmZi0dUiiHvobt33DimQCi4kciPInuuCUx0uMGwsfm5b15gBD8cyatLgVwaFLRBlpgqb/fre
keaxyqvNsKQg+2KrjVoXPxTgcbUAUeRNabTYHQlRHoRRWbaXcZV55mn6cAks9OiUdP/3ENvW+KX8
qfuLEsm8fgYHn9Bhi11JuC4RXZ2N1Zjk15bJu+Khw8zWdW9dcsOY5BQwgeN7Yd+QKDGpMN3BtcFN
k4louNIQ+8TYZPcH9Qz7UttUVgKR6g1ECtMYLwGtzgoU0ch5rd1hItjx2tq+pehmgAclP30VH1jQ
dxpzZN9OCSUg+KZl9VoT85W4tD3AJ5LpmYj31gIWygbqYlsMaLtKmJ2iEpmyyWccal1EWp4PS+iS
Xi/TwgHghCMNObIpqz4AfSmyUxpCzEyhNGMRZ7tvjUb/WgTISplC4Ir07u/DMmIlGoVnCkeiCDJY
t11UXTFoT1Qt3ob3D7DGXSwjw7nuuw/RspIWjpbssHMHsRePlrQuU0J83A8LP27ZpPwt9/nZ264t
3VApYm5Qms/Wof0iqyhJfwnJNeGZb8wfChlYfTYogvkzHxNHD/wbIXmIMkycs5wva+LvM8c0+ZMt
9KU5JzVxreWR0q33Nr/9Oj2AO1ReeY45ZYbhZyI67NddM+GkJJH+pnzU7ebXV4X9HMcP9RYNpX4A
L1LkQWeWArjQSNddxkJBlNWbgs24SqOEvWB/lZnasKhf/wAQAiPhvkTV4Bnk9ZiCuJIVHq1zi5ui
qTHXTKD1QfvpR6uhXSO2+k3zNMJNNyavlsV/YlvNi+8nhqqzSwfnUEcWLyjKuVBi0+PGFF0Nqi6f
Mtcyk5pcjpfcG6fY+dgfAWymPilTWCEl0h5LayEfBBJtIjwDOlq8mCIvwIKpkk397tzJ8WXaLT0q
sDCn6YlUmwhaS0WLB+imoCvpvWFGYZzpwFZHjxou+XuPCj7AExvMFQ8K//PGdRseh8A4A5k27DQ3
w8dFTSshqQDdYn0KMxXUEGvc2DZoTZgaCU/05bzcDLBS0VXRX3375TOkpq6MOzhwiMNnCJMw764U
F4qzlD9llISsYkwAbSkL4YmfMLkWop/gDGS+REp6wEdRLkrES7cFbh5Xfb684wcBRUdcD3vID2th
SzvW8tmp+J8Vuu15x6E2gCUBgW9vlSbalZK7CAcxpTVsVAToZwYjtafDpsebiYgPKqD/dyEEHThj
0knVes+FL4DeL9Ah8H5BYSOZDHdYpg28UrCu14VELeK7XKE+JLRYlsWgy652P5otcmHDFheDHRra
/zZoaHxJvuVZLpi+8cdpo6sMzuMyiQ5N5zyLkyukB/BuOPOzcRt7QqEz43C5Jugaw/KnDlHdAcO1
xF87jb8YaU1GmKquBTn5X5PtmRZlVHYnZQODLXs76c97ax00T9bCrJQnS/tQI/2ZJr8/D3qRtyeP
OMSNVV4Nyp300+2co0C6csKmn3cwE8uSbWotDhKrCGEuVkvlt73ybh5ijudjDXf3bVhfsXIYPCIt
0zcZnl7LQMqwANpt8xduGG5n+bpzd/YIj3s4+ln2uuxyrjaUUUYOKvoCCKV1Z/hehlT1rx/5rMyA
7vHqMxpyYJBpHlHWttpKTsZWkn57OEHygYHw3JT5SMqnO0DOD8NBVgZ+N0sCLMK3IlDXzc7n3NCI
grYN7CRDT/eAhXSwDi73RptzXICdMcEjOigI8YmxzXlGn2uFQT1q7jL9avmoNeH5qCj0ADewdKuf
n7B4Y62LaTe1kTE+KYxAtpLR+oNlIXyAgUuIicx1szUazWrf6OSkMp5Ww+RdAecK5FS/kY9ESjnI
ELty6M3ovWZQMwQhvXoE1emnz8w1ydrYXgq9qfKZ8Ir6gsBldK+xpQhlzwL/CM5IE2Nq1LiO0bkW
9X8iWcBHWkvH7J9cxkAhT9l2R4dIrq1lfJYLPluZwrCeB008YRmqQqotE9Kg/4Li1yom3pUNgnEj
RwwLpb7FjynxdH6A+Ctoc2ZwC4uzigIQazn8NNMePpf/Q9KV0qMT5pPCxW3rdCsW+n5bbG3TnCPg
oX23HKKOZ3ZgEmYVg+pBMP2icrCAWWvuO6DqnImqJyWMjbxN4uLFLZQie7a0nPbxFxColEeVDo6C
mCffRoKifvyLanRq8AxmUts3svPF0dj13nVWhJj3Mcd43Dyw433utnoNGueFPWBrTakAebgaXONi
B/36lWkU7Kd60S6z8VN4LzaVnbQGItsyJm7hZzHUbm7Lp8Egnaasn81qfs9XeJWOpwi/WGJ+UfVA
rWs+vBAQHqVKaMIG7sPA9bSmwKd200IyASTVV1F4BEBURUWnc67IUkS3LqLhzECLsBXragp+8/qe
6w2yj1AfRBUF/kPI4lj82D5W7mrbmeX+HQx8FQZUQuvIjjt/OjOYK8lcy5p1BVQ5hgCsP+3YUMMT
IFBd4Y6eFJ4Ssvyd/xB2Drd3uu8B6Ale13GyH1ozN2v9VrHyDtWW/RZaO7SzAA8Sw4IazMM2QaLl
tehilpDcTQ7FPH8sFLL3/NeqQAOlTeeL92/r7uxcATxXAwjnpTdClz6GOvCP8I6BPJq7SisS3HOT
LBXSbK08cvV7JlWzqsy8P9pMt/rHWasu2XeDbIVFD/p4J9NQp5lss1c/UYNzKXZWCnzFneekjt8B
NPZUun2rny0lvhukZVNauWqx5WIE6E972Rkz9mC5Kgly2kTA4AwSFbp/jfOBH7/dnvObirIeewDh
DvD3Nqfvm6Cs2gXoYAsUVLoWe/Eeqdy2hdSv13MT6Bb3A3yWrQxMzdHZ+6TPmfqWv2diQKm/KbTM
Jq020r6BKqJtdlCp9TMRg3ZFgsGl8D+BokCRvExuhCfTGNeqjHTip2qZ5jJDja+1ITwSMPdMMnor
Mt78d8AHrPtBo0sSe6CciNsoBx0YaUJTp7iV6AdQxRINBYWow4/kxO8Uy5zGePEy9IyEyy4dVdSq
pQaL3K4weT2FWXSGMoOTDn8fqAnBb1AuxUJW3/sCMMXMSffA018CjX05Ogqw7LDTcMCaad0xJkGW
EgTmwypU4T+YlDEAQiA8bRIX7muJUtGKvUQ1kLWgYbhoc68g2WLyKAazQJaGqq5fYC88NupOF9Xr
tHyZDLG+PPpm1q6P36Ie9MUFxK8vhTyeOMcrKjb9XGM/4uBV+m5hqeBq3MytfYjolsrmZt50S9le
caVSJKghRlLnNLrK7Sv0OCC53Hb8l8XQ5/OxE19BwMDsMmgjx4NVl9eDsufc6wxb37MO62IXVza3
/Jh4ccxqycUJORQzmAnd/9sFqvsjZRuK8SYIinWdprv3kCWVc3biLQNzG/lkxzdSS9eTJDyQypL3
sMM/4BtTs829URD6pajK3ZR3pkXB6PbrIjsXCpEaf4BExXUYPFEgsnNDXAVHXL7bAPCphJHnjoYj
+80YxQ3uJsotcYrXEl44Hn+0IONsS0jF1P+tMRGlJ/qL4njXshoz/Gsk9TmwU1tyZ67aB8N/uQvw
byUPazcI+MapdMoswRlVyJfZb1VuImtYXiJlBAMdSxljX3pD6FcEZj8tMcDJEcC2SwYT7ukqjTsc
rGCmSW79O1gnfyfyoIJ4RgnzipdOnK2MeL14NzuGCY2rwe4zrwjrQbZy+Sq4gVLHzK9/CHFEQJ/E
fvmzo9ybU5j2cu3dn/GmsSxqSLo5Po91fRc4U70adGTFHyl0cyGgr1LePTyrR+b6RTO0g/KIj8TC
vQTzPuGXP5mrV16A3o8U3ybEpVBrCVe64FrGt4nvvT230FWc2JfuLfZ4rOFMqV0RXR+r7Jw/T78m
qHQ34TThy2TFWNxW/wXEKBgjBI9j5vqgyfby40ePG/vt3b5bH+5FangaCxeEdwT9IUupyViLi0Ex
2FMB8Udb+F8nVWG8jWHR2gmpjaTHJtUvwzszzSOqeclbtaXsCOynBox/vlL+GfmYBa4j9UnVvpZ1
5VeSfsGo+/DdfpiJh87HYdqGw2lyiCZrLvOt8QzJteytAhdYqQizLWu49+mnTb+HdRLzlcywd2kC
0f+uIbL6M4lJe9MOJcEDLOWcTquJKv725FggzrYdiOe6OW9aA0ZVfYPZbjXWgDvSPZLQrDzKhYiM
Xh8vlbkZEEHOkaOioHjKbLMA3RuIOHY6SCSol4GFcgbAZ28ZeJ/E+LJdjEzgak5juvE1G27O4HYI
x0Zh3rCyICqGYxNEpxKTHiUp6N4kUt4X5U2Ih1F8F/KohGiet0ZB4jtD9pDkmBCkw7zQkiSxhBJV
9YHqrjTUbIVHwo2ytjAtSbUdPMd+fLcwmgYy1lWv6wWOhxXLCbGiL/lpa8GbhwXwNzIZaeBQXgSj
A3SZzFzB1FpfM5/OJHXolQACjMwpwyx91L/nmwNLSgYGUDrVR1nWE8T8v49LDbNLNJI8KaTEia4o
WmMQ7SmJndn9rmeVmPODoKCOfk6fhsDsgv9zpyWaASNSIqPckOR6Fj4B9xtNE/Es2r3UDAeSxfuW
QAu5/uJJnWuWfbZDBxY0mXX8xnH9gG/i4Cqgfp/n26Pmicu0LDQWa0VTNqmRKXN/ORgLg0Y1VkmG
iAHgeLp+gt8i6owGizMjMuxazjvJX96JAIq2aJ+tkWewN9xieh2IF9jqKqBHW8WS+UDitT08BL9R
KAG5vORORsMM3F04LPR67zOWQDKZSw3yOV2rzAyfwQ/KNwa+XK6hKtSUP8o8Ge5NdDX2dd1Uo3vw
Z3lqb4QPIK02Uk6GAGJIEAB4ZoXiJZc0YtMR/sKK/HBYX5UUgQOUDRzadMByu4F+CKMxp0lwDOUl
+L0liAEwG9UQ9l9HcNQz9fvB/qAApUL1r4bVkaqpyCCbhSTZkeVUUGMZ8zFisF57CQgVBhnKBvso
dWNEqWDiKJUbIc/HUCnb+QsjuNaoIIOB0Auvrfq/fp5/3eISTjaddowFbo/tL7teIBs9UOJfAUqI
MtaDWm963xV84iNhtbRp9/XEvijCc8n98PaogBS73/M8u/x73JTRGfi2siCphNI0VA4v9knXcoYz
bK9VUtMBX4fHhNVOSdOrQ6eaRxM6BZkw2YrnqbUsZMT85Abe5AbucNU3SW23Qs148ajxd/Fie1p6
tVxx+vUIXOp+xJKtW8VhyqE6sTL555V9WRBaigX5gocXylygzilhUNPQSEO8gUYGZ59RU9JB5mvy
HF5K/YkcmhCqjUWDQIVr8EOJ5yjJTeYu4ahINOkx15XGJqGurYbqeCMSSMKNdRxjFyNSHvobVFKr
Ij4IUDj5E14GGpOPgA3Ec58M3vslB6W654361L5X4EvOTjlI0FWiv2gZlfVDUmaptogOc1kQyZuL
PSKAfvpS1BlUVBqPP3+NQxeE0Wh04m0BTHpA4AizJ0FybM+07mcVaKC5uCDfcNEflUAubAezsTKf
f9SRht4lkGMp0vON5i+wul35emEFfFKpHL4ZFycgiaRxCZvAi75uGpVGKuxWyw0f5lyPOhUS3rOZ
Ts3iqvrAo0jBTqRMRMFkgANgW23+OzPSHp2y47dhyP6BzPagwygw5ALFIjgaxDmEKmmZAO36QtMa
rWTTstGnmTXXXXvZe2cVvNhqaSYEWMLTDz8yDXrMijlqk0mQUh6NDU8tIcQRsqwdkSg3KbuzeOo9
aK9knIPfbBxFXCSafxXQo34Bm0IM1Ok8iB9KtL+eGWHyAsbdFS1BUoNGQ1+xALQNJclbDLwmnAxg
MxlFarQHOYHWtHnsj4v9IDnrhAUbZq4OToCE4D8ZWH2Ovbn6zw7QyFECGn5FQww9ZvCCtz/QVOcY
9kLUUQ8EVc6PHgtVYhJaF/KZDw3U/Jrg+LEwZQqhWKmAsSbP5aWHRMU73Jw9MtPDEkCK1sfqVy8z
VAaO9c9SjhvTSKAaaLfGv/Yk93VaTGOekGsnVRm80PPkIA2v3kXRL68Us9L4/1AZqHnxx1OrGX2T
B21tNbT62jFAqHAW8uOB7UAARZ1phyDdcBthKJrpK21cEnxRrzhHBEehTeT7SD9r49ZQhpah9VsJ
DtS3wM7H4h3ZIkN36EfkptvkP2peGnTkAuV4Db0MclTta3+3Nb5+L3AWAeNB30hLn3skTJ6PTmkI
c7zsUg9fRIOu9tzPsweG5wiVjpTgKAcfa4El1BHAEFjepXdkIA18XScepWRsOPF6d/tao6pycvIL
ImJTtK3exxVJ92kGj29Es/B3+byz43Wxo46ka6VDvI3cCqmkGZSVH2Kk2xzsSoTzF5deERvvXmSW
uQ0XiUYqbsXJpoQD/smZht5ZrkHlIw7tMptuSgapqQ6LlDjkexIcUSBfv5iA5jCsayQipqAJQAfv
r+IARVXYWhjp8GuTbaIMjKTxK+P718tX14wJAM2WeukPTJeKFgRCQr7y+Y0mQcNg04tGkeTquuGN
jmspBExHNgE+hwHNhO0UkJRiHhi+dqZHSGMS7oGlLAbBqN2QbhoznWtYFc54Z8xX218D9aekilBW
EDnD1PzDfMF4l2asOX2DCw3p7DbJFda6AP71gWxmHxKxzlTPHOePjLE9x4sSvt4xs1ic3C8qkIrk
oT/wVvPbpuJgY0l4Ku3DQDUN+vMIBVf5+rmcHvMtLj3WpbaQijxS2HZIiHWVOteZYhCUA7TB1BIr
IXTS6Y03mEJrhs4JXbGvBDFYLIsK1Yk6LIbLA8ZpOcY7XZ9D90RcT5oOX1pI2ZEdU1XsMPIa5bZS
j6ZIfgE4XL6j5l37V7BVnVWBO96+wnqoVRr3tzFqSXLTQu/HP7LrAwxpZxWiqzMCwIYk7v6pm7gM
LRFvGDYjdGePymbU3q5dSpQmkusQiD1gJXCk398e6f3MSa5YvByz16c9GfMoAwooc8VwT3oBVbYG
IMc2DxLfd5/1I6Wr5t9IPd4jgU6zX14923oup6XOp4w+eQh+2AWslOcv1YvFxw5o1eehtv4/2+Bm
83uhEsPhBK6qZAoLROZHXIB6E59WNT79IjlM8zZ8NvWVTdSUFu2HlbxUsh1nklO8RcbwFdk1cz9+
TxY4E4D5yFl1En+l/LuQa46Hftoa+7jQNimxhue2rNDwUxgVg44vYrU8Itj1cqTGb8UxAq9RlN6s
ywRbFCRdFRDUVoH9WAfqBD5Gunxvriq8FYJb6a6jIeovC2R5PePjlFMadgjK4I8oB8SfXoyJRDdd
dEbyz+skrfK6FEuFjbmN2gGI907gtB3N793EmPVAbnbRDgbfSi8sn2nauGQ2EHk9hKPWyHPivBf3
V12tRAN8T4ilblGe6ey5Ma2ZDjz9uppu7oRH0V9AdVHoahlEjblbNpfzMkQPoGh8HcG8CA5F6otD
km+nqi7RfC/JWbWVrubAPuQn7Hs7rghU9liMfvAjJwhCnH2743lluIZsF5mZo44Ihi9ZXwRc7guv
SLAeSnseUpoFXGjeZCIpeLJoxvpqJYjQBeOSEZCmzvX+30vApxwgt4gxSFq19znb/83eO5DKUJBc
Jr9f2dwU53mdBcp71rR8pBWo9cNKXMeFWjQjVpNtmaVBnizgPcfomPSNGpal/5cjgpzQDSNspBG7
/84jfOlzYB/B8r+ay61SfuaVOGGuQ4ERUKasrXqyjuUOhzN+4ULZUlnihAXg4DDE37dV9vQl6xxj
lFg1RKHJS9YlsIRZ9bP+vCayTz6xVi4h0gHXkpfrVzk3wtmWFiTZW4KGeTXiFh1NqKYSMJSuTM7i
QDGshHrY93YZz1b/SR342BpAoFoQtsLNBD8N+rBR91o3X3whjV0Tcd/YV6//bLT5fganRZIfJVr1
uG4KTx+Y+f2o9xKFyB9EvM7zct7ajEhV4B3R2tSGnDjpvOx9RHzOmVqGD6G/WBc2O204mGEFlAPX
FMvSrbqiKgf07d4Bl4dwooGzDYxSMRZdTQw2VX+rHjRm21gzCMoQG1I3SznywN9H0dGexc8VX1x9
aNsUA2b7NYMvGkpMdxJ9pw3P7gbVYyJsNRUC2Fn1kIJSLhrVAxXlM+MdEm+HS9GiEwH6BrQDltj7
4kDi5TqG1g1swlTniyE9P4+3JysCTD7OI160NRcxKdC0cbNIaQ4mpi4SiFA0HxbN7euUYb5srfOp
AbOw9nExKkGI7iwpmQEOiEaOL4FnmPX2jmsurZwrPCYmM0UZwGatT4bSpO1E2SXtfufomc1AR2dZ
rfWGJK/G3nhXXAHPmcogGobVH81XpQkOiS0Kz3UVhQt/Zr2SjA/rHKo97Q4qGlm27/fAbAMDzRkA
hBvrPrgDNL21IEDEf064sC74P4WHrgiVfotm2qMP1qb+ya1usYP2sI35tCQdxShNHE7XOfJwYsnf
aXYn05LwjXOKrsZnbGhpWBaz/lEBvIV1EH43tS+0zIf+iMrlN7JE67NnM5bQetWWsJ6BvzhS22Em
ghRrcxWw+leMSBvcbx2u0PFeK0Lj1v9izTMGx8cYgOMc6mEq+pQ1kVmFFVFpheCWHYEk1Yjw9yA2
oZOrUBW5qHP35C5YBHBU/6fe9iyV2tv2GDWGkJu94XSuXWTgNKzsjRIvHH/23WWbEDNucoZsRtIp
ujXDepDK67k41Y+6LcZddWJYadradR9zzx/pBhvy1vWoe7C0CGIwpms8Edpkk7a4MQKW4ibjJu0o
WEqVWLauqduv/aWW5j+Z8feI5AWYU3/15kl6m3s+fLuLqb29O9UQLrVoczxHloZQHolE/xqH1u+d
ifHnbBIjmNIAm2p9Jxw3j7tKSqd9TvPOVLq5Hv0skmB0smhCITxeKcOv+5aJZiULzyi/1lVJGm9x
jmWqr1co/ez6Nyed7CC4Xz8npLKiTduHb00jAHO1RS7larUHRe20GJ0iPRMWsHhZ13yil3ardt+Q
MEBJm8QKV3qAtFlshtGYqeekxUjQISI2CwW9gyCi29EHiuNZ3+jd0a9Ra4sHIUMyCeUmBIOlPFPy
myUF2lC/EhrsUdyKY7/P8wHp3Slk4/+M+ew8Wqgub5m0XHxzum5L0JFTzI3gP+jGHYySa7EpXHJd
SWGRfgDsQePOJaHmtGARMjkDIGbGkgtSwDU+5lOoUIzKrm+HYDIdwBP1mvtb76ZBoZfIkvQEI+O5
YiczYO+Ci6dgihHh9wiWhAX6nf/ZFc0JwmrHxZ40URNrzb2fPJ3FXswFo/snp4nMMyPQ3gB+XVcZ
anzqimH3jyAX/5BZNZ6DratVYHeJCgygSk3aSWg0yB053SuSORA4g9c6CMQCGoNZgJjFwRsUaC3b
ynAgUF52wBIPmWa3UnlJ7bY+j4D98GWvSNOkau4vU0ocB0/uYN93ydOsdqqbm2FAXdln2CxwFu9a
Rv8/yH1o7kIRbie6B0l4ZHlm0sY3laPIjN6xtMg35gO68EQlAH8Z9Pq673idWS/gqgXsqcGnhiMG
ck42HI03yy4QlV3Iy+SuHinNg2js4YPikRLuoJK7JvDnq3vYHczDg13tAcMvq7mxYb241kIsmhr8
YPX8McdW4U+DeiXMgfsz+Ix+0q1Cj09IuIipjbhl4L9DDSbK3tXWsbiuGwoWdjDgYe6JC5i+XlX+
AMibRac6Ohg8u50+5klpk/6jdtgvuae6QHMi6ITnde5joKj9RbNNzOijl6c6Kep29W53zNYERk3a
GK25X7NUrA8fh4mj7owc5qMc47uUYPdGmAt72DgzNrHV9Gll9tMtKTQxY6GnRdnhj/z8Lq5iWGDx
1L1ZZFZM8jJTAlAkXZQNtJgJ45svkzBU2HurpdloV+bWbeLUo+Y3Idaw7N9zi/zQBuXeNL6DhOcZ
7dJRUlD8Nroj5JHnA55G6aBT7qMUdw0vDZ6rjPesWUT8WAsO5r0GNgvnDsXSRkHorCxKYwC2qAt2
vPN8w01QK1Zkc9yb48dn+u99ilxtARv9CvbFqbDZm0silV3vFP+0wv3x4UzUWldScfvptNbZXlMq
GuuYxMqM+3iXRc1NGnZd4o//LYyPw2ANcVWREu5EuoaKG/wLb8RXFEXwSlKebMecO2ZC7wuKUD1k
YrgW/XZsYJfkjccFnr2CbiFMu5kYYqt4CgPGziTu+SRPOKXwGEmNnmZMNHnp9AC02VnCQm91Wag1
Z/UpGIita/NrEkaQXQTXb0Ip8qYKx3Qk6sESDPgFiAX3JvgphyVuWmCD3dzAyhqtz2d9rzzweXYs
VgwmvmzqktmepNZ/YCCRMZ44h6k2Pz1ToyK6jncm5Ov4CD4Ijcxgwo5Kn76sxSVPU5e/V2p+uWxv
XQLw64QzsijtaL3fP3T/VMXJAwJhLuq6xTQ7/TnB+dwsk9kdt4GdJepUFPyc6BaBDspURdZy/Axp
cBYHbjIOkiT9K/JSRS+pqCDKfNWzvWCwNIfb08L5icnoFtMYspnIrQU9pv1Kvfp+JPXlKtLZHU75
LE40MBV3Ltsb9KxPYls43O53S+oCa7eK4485G7VkRFV2pWYXUVBTuEAiS0GLLr5LUfTW57IllQwH
nJbNU6rRAsdV+9qs33OfbidKNWVYzebwq4VpNTBWF9t6qYHOSWYf3TeXQzRm5h9CDdmmLhI8vCPL
ApaUkdgcznyfOHQVw5s9NtX2FNBXz3lcFYMXsRc7+nK9XI0xXUeRbDkhSjPLKfG7E8fGGGMXsBDi
bOnu8jT9SL9197wLl/Iwh5pRrsDKTzL7tQ+fLh4ocaZkrjtxl6dQqfkfbE3zTeC9bkMMdx8bpjRd
o1KP4C5/dimt4tS1U6apuq7upUFdsk7rjShZZrUSP0KCiF3AD8Km7sqOx8Rhr6giXIpDKGJJs9xO
O+JtpSk2WL1D4A51tGlzF9KtYXxCF/lw8d8gTmGFBk0xvVXyP+0pb56y9fhSnX1VpTRZID1sopCj
6ozYNFkXb8Oix5r63vd4xUv4D8ub8qoaIutCM87MfTCi8pW+2iiVZ7fKH7vLVqHO07rwAU7KcEqz
LZt6/yKj0SI7gCVuvGw/uDiqbBfDxO6bihO6f5lle270+bnabELlgAS1espPozLUzd16Ot+QTRTx
Be6ZuY9vyVqMXnFPoERSKWrbfvbAfOIjJMvw7iplmaqrluJU+GBS7sL6qoNUmvGsM5lioPBkyw6S
ToXnnemhTp1ZgIZzloTjqeOybYDSyPD1Aldb/ucb8sVU4DQSTF3U0XyWqAPkeLDGOaDzIilBpdWf
KRw8KBkwmFl8YM7O5Rp5X8rOgsxQMWge5fWNWxGJFAaFKHiX1NCGjYUp5960u4oQb3yCQntmPPzT
avQkavqf5RTQ8pn9HxK4f8SzZTO23BNs4QwSH77eBpvWX4xyCJlmvH2bbIu3RZOlMbW/n2Ash9m7
Hn232x4yTTT2/KBk9nwfq6SEUfd0ZrgaMNWAYefGTjCkasX2v767P28KOgJuCggvgHSiwT40LEIl
FYwJXcE19nWaJxi+4+6k0eLpAsPiNsz9fd8V2BYtdn4jT7iatXXGqbkIj+QmO2He69zZn7MWCkg+
Ot+BQwqpxyGBODXx8vksdTpTEI2ZocEfii3l3rjjlwWzV0KFWNtFzysyZDOZQJEwl7F5dUnjBU5v
sPT0K9MOMyBqc/0Lvr1FBgsZlObBI3nMBnhZIjCDAYTgiS1X7Z77zEz3IV8uaDTlaVcEPWWIEdhB
unXcsxqy3XtWDyuZERMjrPakp1Cqcp47gB9AWsXf0pUP52k2rJ41yY9kRL8NLpab8arM42239Try
AEa82jQ1O0saVatNcE6CL6e7+p+SA8szJkWjIH+iblGO7CunPZLK1hxl/oqnDirnP/oHguz5w2At
ybecjq+wTbs1xVd013ZDxFQjAlAkZMwytiBsrS7QIT+Z/xIx4zGgxDx+b04BNgSRbCPoVUCfjckF
5r7jzNG3vRevYtPKnIUuTKSWj5OViUP//SQ0Zjd6sJoZyvsbSL38QLhmpiWAlsPTtmOsYdz4DtVt
CyvDv5+VwcWGs01DR/8AOAmchY5E/qnvntOfyIGkNYVZkaI/6R03KoiYBHQA1OASiB6QzLZnM58E
Pywb6PkPkUsMy3eqfKkirREmHOa/VoV/saa7wrDB5kTZvNbHT5JZWUIRPv2wIcEruxAhWvyNNSs+
ri3qjXmaBzeDOhthz+Z0L0S+vGQCDobpLZbI/vVTf6lZlov5l7Gr2OTLLpZNg2bi3W1oThFirSVj
1lLS+urli54BPKCsJhB/VOyuN2BDpcor2owxqUNujei04t802/OtRjStu7r5g6m+M2gRTG+/54YH
bcDNUfTuUZe9ifqszXiHJZu4RjeZRBGZpLf2RRWXC7EywzzV9V0CtCJu24DHrFZFvjI1TkIXXKln
CMmYY2XzSi1CQWlEjy+neNerIeJWi19va4ye7fH0vpf2Rkdssfb8zP+5qdSfNxq2MPjckBBHz4LW
cs7ZBOzC6h1fNyjwkQyPuTh424NQd39YlSXFda1jTLFeb4SxrWv45vRLPiCf4mZUjCswzkmw+OCX
otVjTtI9/ZrVZVVP5Wq9UrfyU7L/du3rH0/rB+xth6xeFtVqK0l8fkiFlPNI+XT7Z0LpWnQo/FNf
D5AlCzalOogLj/Rcvb2CvozM2o7szZNNIOWFzV742yHYwidkAKoGJHimhVKqeb1GdA7oWFcRjvu2
RFI/sj1pQolG0rZHy7nOX26lQQpH9q8cjID0knFN8DHIYQ+cCQH5c07/PGmv0So682jzZ6BfGqVp
uq81chB629a5yWcVNJnONx22lM64bfMPFB6MtQ21h9O+wM0FTkttqfnazPnB9xUlAw+yjqc0qkLO
HY1XjSCVPtE/ri6stAevO2g4PlQ5AW5El6bhczDO9H8ZSJ4mTSEWYWyj5IAGCioxd/A5QUZ2ogq3
gdDGdICxAX+qeoZYp+F8OXmbljhYOZiIwRHOtPaDpmkCiulimS3/L/tS6wloCLk9+wGJpzWT1pHD
g27kP3WB2IXJa+5vhprUbvjoKsLhZp7yBa17RT5H1MnTZGL4ibtgspaiCEuxFLVfbgDYLz24DZ4m
GMbx9smz9ZMqilKhtAoeryS0DbLHl+brGNA2/O4PvbE7+6VFwj9eJrA0kJwWyHw6QMW2zj7D930K
6hGoklD2YZb2m62hsWwMZ9lj8/XAy44CR4DGD3SHEu705OJFLLiqNTkJysmBLmcrZOtK6D7fhbXK
alad/GfjlBYKkSVpQr7bvJYiNWmY2SsF7y4iP+UTrae3+2qPN4ZSxJ9FJWjn+biexcOuCnXuLomq
/mNaWtQcMrrXex/pZ5Aj8Bvyn5D9B4KCZATfXHbBw3qFWV7TwofGrWaHg4xpdHKx46RGxsPMrwN1
p1CvZ8rfQtbsJJXkWItgjcLr+2xtTUstR4S2ST96iXGjDT4JBycjxhvU+YXBUqJjB0B+E2u6Ew01
aCJjRQ3Yg2Mk71sXzVMKhk+2s3VZF+3t8lu9bq1aDBySIPm746SlKr+iqvPZaPFm8OB7k9fvSY82
daQSZj27MIx1qiGSvGggHGOgByYY0nqWUSVfwi5CHVgWD0d0gRSOOy3RPn6SHM3met9QL4j5LRhA
BgTB3w0Bvg2Z5Ao38QIhIaopHB2cjEbitP2lsJfCfWN9SSSHX9QVNgb4bDtAlr6vNUa75CzrAktV
ypYW138KsrR52T2OqSqp6cH8/f5CvetuvCVS04E7THd1SbWh92YZfu1/gSp76iFJ/XE2v7/5xTRL
M5k8jUYDtEbbQOzvKiSRKdEIdQl91iZmv3/UJfKnciDJgId/Q1bKce0p8mHOXNg+kTkhQXqKfMjc
85K925v7RfB1VQUIlo8GxP5us4jqPPUZZAXAEu5m5gaXiPwTQoWP1vCO6pTdsYtSdLzwW2W3Fm9u
d0s6/kayGvNrO9XhbhszvdTvlgYyZ/T28478kUzq86LFwToTrHZUmbn/sBueTqWAAkZvLyVtRUdo
EtzjlRFlVtgUUfMQEObpB/BibBu+Zl3wiNxMtnbwuZWL5MkVFiQstIzBhL57a9Jpdhgz3snirvVc
DfmL5NuqmJbe8gp+V0D0XgCTdzJ8mCVgSBnV9YlhRxma9cUaYmxAdbju9vD1yb86V4xgf1ksFUSL
N4PcU/IVOpVSQA6ZQZI+5522Ju50X+V36lm7LZhFaYEM49TQSHH1yniO+wpfMYS7zw3aLmN81ECz
MI5jmpY0eB+wo6xfnLu3eqm+KjCS+BVdm4+1wMrEdxx4NBQPsMcZCTptGF/jOA57qO+11yLLjoFL
9d5PohaySsOElXsntCqY2j2oh42W/c6hP437hWt6JFaC+cCdPvXeG5p1P2405jAwWnWS7kDtRHFJ
zU5Zm1mP44/cxt70XLuE41syVOc8xTFDbDiYQAuTt6OZN/5/7WpxJZfcoa1IOw6il+C+7dEWvsv/
RD6yjIVUJkAzgO+fY1sY7ZgFan9EuUm/+wrwDfWELiOr2sGx04iCPUGfXMehC2CTbdHl2poiRxsS
3Cz8wubWPm8OhVn3L7ncKHLmmZCjZC05m3QOuFf+L8a+aNmSa2Nox4idJVBuQdXrzbMt9VmYmIc9
peQhZsDxPGtN4X1xm1wbi+PP3pBoPxN2BsKchpEPT2Fwnh9KqQwPMK22fuG4txplIKNcpldIMBL9
i68lN3Dzpno4JMr2vILUWn2Rz1xK4OB7wMNETCQPAi8TVXxssqwSqLvMpZkJDPn//54gTv7+v0Tc
R7z6qs7NCGaUl0iwviuJw5BIM8tgzUSD+DB7nX22CzqX3YYJgC3qpAIUOTrIf/tTKmFoJ2iP9nUl
LutILtWol6vYGTreq9n2fWn4/hAbpDhkpHaCWDD9fy3Wn7xfSWFaaXQpZGzAAaTf8nLWQTN14ySe
tdx78G0RxxoVeFrcGDA7j7H/afTuLsLPQGtVevG9OU2y+X6jqvQDqAo0AEn1TXntNmtOvsPczXM3
8E7QBhgjhW9Jnz1MxDolqkpnbd5VumNxMebCdonDqFoKWSdOTry2L6zPfwG6/FCQINpSUohMBmqV
KpzttcR+O2hQCEqT5ppCkKtHUkHQAX25Zbl/M32G6Ds0b5b5/rBu/E/zVfznYnl1cKw8icR1iBaw
OEmZBKa6bnk9jsQ4wqAoYHBTuBTeNq1NJUMAQjQi/oUGjmDkno0mvp0qh+bLHiKhcQQq8xeQ39pg
7qKNSB6Aia11B2rSJiaHqoMpARRaF95MizgW8sqFR9Ooot9KR2Kyrdk0ebPAov/FWuNzoxWCaMeB
sykl5VwGeRXIueSxS1SQChOw6Owo2YC81mdnNPtijCbvWeCN2ifAOv2hJJWQBSDPzyJX8O/O+BGZ
7fktS7KkajgVkncuBeqEiy/7aZ4Nxbn1jga5KfJxP2e/dXDB06ld/RJfJoYA6QeG49FB9Dl9qav8
pP/Iriwu/KNw4OqWwE2Gb/64pazl2Q2anjYpFVfpSD6+bzAvI4iHncdLnb9zQZqEyNqCljJZkDu8
uZhz5UYXZzZupF6T3elX+VFZ869+59oHs30eRuMHYX+CTYXogsDaRCsywjSVBK4Bvam6NPwglXyN
DI2qstmdy/UYQCHs36lf1b6MyfSgVp3d/G7hRN8ujN+aGhUktMJtgQXrfIl2Fs17DubUuYetlU0V
1Tg3/iqSqsI0HKT7Nb/TsPcwi0+r+AMnAJeZmlpEWTUSbeYxahXQli7JOaZ+boahng0B/RJxGQdL
YknYrwtVInchHub2wCfCGhImrihiSGfcv0j3ekyVjQhPumoj5Yp2hnu5cqDzoGwE6qMArdVftvZq
jBnY9np89+O7RYwjmm2pRHqglzZcC0vdsXElXQ9zWpvloCLti0MRhz6QqqeKXzWLishxo11Fl2VU
2CQ/V/gSwuTqdQVprfiemrDjrD5c0QpYxk6eDtIXUktIgBGdxJT5FBSaAb37rHJyPsMLQUnreQRW
EPxdNoO7SHh7lEWd0r1JpY7CDJXKqls2yTFkOGEErBS8UV8ynpjziydvFh+DaR//DwTQT0h5SLMY
v4LYPlIAF1rvtsQFj7EHPVws0U1ZU6d1cMuzFKrg33NgjSmxBVPRQTcZajE1A2UynnUYof3wPoQI
fxpPshj1y4hrQ5NZuDijae3h0PdNZkmhH7WV8no5nqNYab8Obmj/qySJhJ8sDPfB6S+RQML0WWnu
ShNwYbCKxQbnwTp8EyX68xE2efyunNo5aK9hiy+SLI5w96TP2eHbDLYOHBgkT1q246G4Kt/BpPkK
c4SCgwqVQ5g2JlEYjFS1eB6DvY9xGEQPl0hzYN4uAPL7ikJosqji7dfjKgVkyfLDWcEuPYAU0gFr
/9KdSYVpI/icW6JSGcU8aa/5HqUmAMl04fuUx0p7+cGGetzerlgzrnMUiEOMxjAkSe9xR/ZFcOYO
S5apIukUotQZYOnHAa/ubLkvkLYKHaspisESUEDTZ3O0Aw4LAdkFx6IJHSf5Y5x1lVWfiRj69qnj
+ERj4es9HlD0Ky1yctbygEu8Ptb7Vdv2M3erqdfkIS+hV03f2Opd0QXhmKcKtaQ6ogIwDIxdeFLN
I1iAzUxsvuWEzxDOctN6GWvkuD19fJO8qDIi33oI2Y5dR2JlMvbX1c0OtqT9bBE6P9/hffDZQXzR
voJ/AhoJQGYa2KCTgSnr6RZRQ8OrTiOBwoQ/wRkw22aa37N+OcRxXDMdarRMNSG71xp3Anl0l8n0
tuFcesZmN3+lnnn5dOiYuSc5rc9txYwR1+gx4MAMDpgCjR4t70vabFsOgqJROUpCh7u8Fr/Nt9BV
UWLwB5l7SjTfx/YzX5ZmbjHqYXwnXRjW5PhaGRb3EYhJ8lOCGyDCdveEfF+HRbSszg4PuoX2JWbj
67875rQzp2Cc3l7aviVxMsCjPeK7efWsdFrfRciiq6RwdUeZl2lfVWt/mJeIUW5+ed2fL9NjpOHU
1/dKaG43s+HLpx53WoZNjuMLtS3R5qTb5ecBl2nWCfXd5j7pywGoEgVeZ6Xypm/SHKuVU3HfakoQ
RKPb5r7w89VVBXb4eQMM73Qyxij8nS6yFk/locQ/XtPFeQ5W5jYZz5AOU54zHyIUyLi0KN4mtZ7j
aq6I14bbLsD+ibbLWcnJX3v1hwK7HyHRUKz3ZkiYGXYR9eKq/9yHuPD0bUiOWAc8taZVsUt4bKEu
9lsCwlZEUxm+qByOtyQ6dkdLs3kPPCD3WJIASir2TBeuDF8AqLHtES9oBqAxCGIHLev7q+i5yF3h
lbpYZe0Fwh42Iqc5LeACghVLHNVBA0Io24LpRwtwMsdvL00slKipNTpyJ4g+7SOlJPHk4231EYkf
Oog4o80U8IlJ3wuN98f2lo9GVG89xFvn6KDdVMwizcT2p3m1fk/fVN9ATu1isDfwB9o8LnifVG7d
BMBw43uYy6nVYDIrYN3RUWuP0tnJ+Iz92Zy1myWF5bNH+rQuvV3DKiVJJiVMBmZlDNSPZ0vMcq1E
YBEpTDKSBSJ66+9v1qSyVhMC0EdAUhwHym5bO5MWZQqEGTOKKsA8VS/37wxKk/RLMmiu4hphb4cl
xBqj96awvOF85llltIo/DGeIqacqBJiN1Wn5EIrY+ozvq/8vOBmHBYf3l5CLNqznQp9rzYqQ0lY+
cK4or6mR3pn5vQx5xJF07tIsWjhAdj5jFoc8nkM6vrt8ok8o53CFRczTS0wvniqmEWQ55RH9qQs/
9m8x1L4oCP7JME2LgMoO1MJE6yzWk/TM6VYNAzdHw+MOuUrrPhH/xsj5Q7oHlTXEKb5hzwXTVmbE
RRGQLmgLP+lEgMht8hbl0u8K2DNxqopaB0TE8IDl7U5jMLRO0LQ00DEIFC+jab+r+B5oHXATlcuf
KvuFSzcW59dw9f7Aab97G6LA7EPc+cFX/B+mry43Q2VtwXmBsJXDRk8uT0LNtSpU4p/FS800PK+9
LAADE5U0xtvBuzhvf+QJ4WDrTUvMZAiRuOALSwn3fvYiymHVmu2+zLskfPD6nMzNf3OWkT6pVUlp
Odb9qWZXe+v3Yxo/x2Gb+Jkis+tgqa15Ttb3j3RIleneAz20USahhPXkVgb0dFAPuhc3SYWuBwTT
bnTB+8lvAwfnsurHy4xhX7fd4wOZfIjkRCA7HZ43eOchWVFwP+FNNSkpqFwKZ4mZ+3DXRIeQDUzS
2jxij8xdLIiN2cqvQItIaFcww4HRP4LGFDD3EjkbGxijMW+YJkdPqGbhn886QQ2JoNZ0aa4z1HaC
B+RocolSIwvmqRNXvEnrgdZdYc6zLK+7xhuSPmFbSBWk3H4batW4P95R3FBk7B9XU0gxVfF/IWcI
EuX+xLICHsz6V8kYZQhRa89BqeIFsgeiAQOojwcWPp1rOS9YBO9nhnvWH13LSd12TTwy0kLBfLdB
xSlK3AfTQsjbJ1yJPDzjqV2Hvx2rq91ZWeCxi9QHvm8OFLjZVzI3BeC1oV5sNu8ZDcPqZTaEXYo3
zoth11wr/OVW6RF6DIXX+u3t+jFOIPt4ZbFk40AxRVvg19PefkVctHUFPyoheO1RODjFaM81Kmje
ttuS/oHBEohxyO3s4HPI/nOeaWjNt6Su+c4Y/zsnWoBjYQfCFcbq3fQ7+AraqCnvu5r/YyerEP6j
RoV/9xEPmUjtUfnlrq0Ao6igAXrz8fcl+aEMds3bnhbIPwfkPgnZjp2x/YvMh+d0AM62SvREZS+g
YoOvXFuYbmsiZMe0GOw9vi6VIgcZR4XXWA8aCpD5hGpxBJiYAlYjToFu7CuSX4W2+tQ6d/5YMMrA
IvywdiDVnlZguaq02pM8SMmkoMPpc0QbRj2DZetvZj/iFYTfZCE9q05qvTYGusPfczFXseuC2JLr
SnvWPeHN0vXlPw/1x/w44u5eJ1RCnffYVfBn9bPHK8bE1fZq8audm29a3it+wCiIa5BU7jVAaYLg
hzNq1V6qACfAbiGemFqN8MTf+uOeghbDhiEvvgHHFcYBHB6J7UwEFKkbay2SAjlb31C/UwTQwh//
OnhBi37N8cv4U9MNj4vi+9aIBoRVcIkLiEa2JWIfll4VhFGGu0f/Ia+G3dn0RYLT8dad7NzBHGVC
mzYiERiVTPBK7JR/0coHDrGaNkEeE0J4g5J/tn5heTHF7uanTLp1J+NKXfdAryYhnnGs80GD037s
hDcVlsiCAcg+fLcKZA94Sczz2dup8aTNqHgNR+U2KkQeIC/7olk/GDoBkwz2P1YenDjyCLFCrtMC
AFhkvEXfM9p6jjEkTIkVfCVNXiyHtGhjarXK4jtAd4Qgb5UxIsNINp2WbvA/NtDgmrphugGsrzKz
BFU06jKoh/DfHGtiay52rgFKZ2PXOc4tGdWVcaqtG+mU7g5uTaJkVDFgKQUFyA/vA0CavEmhhLUZ
uwYFQ0rkaRqiodbd5Nwfa0KDkbXur/fMx0Sj8+FEFzvonQI0iKwrnyIWS2mS2EjYaI/IdbrgZtMY
JiRmuI4OhZF5sm9bhYokC48RvBGhAuplhEzva5CZx5e/iXqA/b7kiaMJDhpHUN/oNp4HfnG5BCOG
bd5MA0bnG8h75cgXk72z6EeY5shBt0/RjmzYI7izbhPvIHSWNsshv6R5qirJwzteA32iOEEBDngG
szfAHUtGhugfKkZ0mz75cJikvwR72e/cCp48ZTvNhKqnzNItjLzJCp770++18+Bm/gCS0zhpUQDq
bTHB0wAd9Bvnao3b8OtxcLPPTRtD8euch8hX/Qwtz424dt2zsxeqWeXxnlSxkAA8AHFyCg7N7Rlm
jqyvQ906uLjd1CDJJnmE3IxiLGAMHvhtR2ipOBPipXAWm/S30bv6vM6rAOShFWEEMwjVa1mwQITA
9N2eivxyqvSMR+nJ/PjNm6tZEDTywm5Hglm1putF553HAc9tgIiINfTr6flbaRd8CjAeoz2D1yGB
npPRI9CLDR6llNSw8qa3NuVclOdFR0j5JBqYy6UpYCrs0OQrp7wzqtXht+uaPEHs46+83ITGBylz
KqTvaazCGX3ttzUCqV364xBOIv9XhYqKKOi9E9t4wRH2BkAJSZcCpuR1oECpOuQPeh6HnLL0PiXd
s+xq491PAcupRhUt7y+Mn2jGApBmyGlhBkpkARXWdm5WdzwGw0QhPBf7fPIeggigBuvkqpLN5P2M
w1nkJNSUHudhIk6+GVEqH8J4EXKoWQ/botKiuZIbXYKbFpW52MUR5rcKx6Su0jD1+aPWR1MVMDeo
Koe8DEBDfKILu5ywXPecLROSPWPOoXRm8kQ3u2AfMiu2ZENi/f1WUX7nIv0tMHDtuLBQV7dA6AB5
35+j4kH5qr6hR5Izilboz6rCQd7mhDgEUW9HKX3PXEcAexp8OInZAyu0MzsKTURgjGnxNTggauA0
UODXDS057hMrRns6CBcsxP0V5D0RxlpzPPtZUhnZa/qTKwCESAkcsAfx4mjxNMhnLVC6jJ5oDtT8
Wa2G5OvyG1fYbtGEyiJre08zjNGg8nQ+HL/007Fnx1bm4/0b6Ey03MyPBwxI4N8M1IOXDInrMUI3
D9S4t4zug9oFpfdUKnxwWrLTZHZmwFFZiT3Y6wz6HkGOjYYgc6IGNPl4bgSFVqVTsoWroVAATuOl
BtsK1FAQOK/uqNHdPo2Vf1gxXDf7KTU6ZH88yINkJWLxcMj91EmCBqyxSKn3TP7BjCuFidaEgWPs
hxRIGWqTHk8UVGQgTKE+K0S6N8eIgjGbxg4Wrue5TRgIb/ysVxe5+25+hGXgFHj2CmISeYngx4id
m2LDq9+B60KODOaEPeldXOZfh7wrEzX0gUAw4Aci6yBQ/PfvVCvqW90bZK1nufBjpZfdcIgfNfbH
YDIOk8licWWFE82GbVCDCE8O4YG7lewWUWyl93/Dx0Bi6oDt++iU9pyrP/ZiJIGEpFBPY8CIRQJZ
FWiwtrkOAylMwri4RMRE6ka6STBjUIb9TCHuqzscUleE27PJRY6FubHHLhmTU1wjZ8/y0fCF60Ob
xo7XlzP2pWQsl862lbpXU8bgDg0XvsFDMoj+yNnr1AgIuxEp/eh/hzs3fKhmpCFhGVTVbW1GfMHm
kbiAzlRkWq3gcFnwjI8w1Gq9lyvXjx+3wSkauuE83OLB3BvDDSA0eC3mLkEew13UPGQMSi49V/Zq
v0VvbFdIq6SB8Hk+bYxmY93LIYozBWnIHpiWOO+EvjhHO95CJj60xEGlgaGt8siF/+/gXBPfCGM2
Ud//+pvJ3bNscXjBEyqem2YMQT5JxPosPzAtMXTO1HpVQzLNWEcPcvriRJLKsuooxVuKV8fFpNUw
gjwUGPHCKRrLebvPBPKtw2hKOzA+5e4Lpna59MAQ8Z/aRnDXtVBDpG64xQbsFPCYNSTOi1/Fph6J
btSmffimaeRMPJfPOOxKy6MXQl9BQ/m4UBAKuwbbuz/z3/b9UzDageB60rOG0BAz/smv97fvsu0u
4MSrgBHuEUBTLzoSj6sjEYuR/2a8H3pd31D1N8di98T/G7opHTlxjaRsxra7GrWAJb9xWXgRobsB
u+3dljhRIwBzeD9UGh7pmkLVwZE+39Y+y2M2FHJJE/DUszc3AOxV1cejBqhJkDUdR8dCwFW8NQKY
BCXzr91P7DdJF4mqKSyCoansZ2d/hs2jc6hViLxyFIvpUeM1DHVyAjzeSdBYpo5+x2bnhkqbt8EF
2yQ5uoiYpdQSlJltB9Ri5mqsW+KxTFI+roon/UocpFv+XCbEIUJ+LS6E4CpymCqUdHhVC65Z/F2C
Oo5dlFU0jwlX+B79l81FwaNaDuHOVMkFPDp6MUuFiexktN/74lgEAoMPN8SJqCgv8l/ap4WZV/P2
LqQGh+DaVNasoOX7p85ygrI1wP2fB4EJSQtquwtGtcmtMZYpu9z2AUl0xC3m0oksqZnudifdqgrQ
X8TNxCalamrT46fTfPiVWuSTRz8aeH6w1vfAh8gZ+KoyIJup8KUAlWiI3vMTomU0GEPHYbRXTlfx
FssSGBeebMVyFhX9byHvCAMVIDBOH/OT4oywbFJl6wMvLgVgX5mYgD7AbsRcUczIlj4RLK0eTIkM
wDrJBZfdkEjTetdb1BLjZ0BWbbS0aTUjuicvJGy3fnEh0ixT0W6EKVAMtjROO0nxmKhrl3UhwL8i
CaUWkuIyKGY/WtXC7kzdib5ABQnipZ2/+ek47nafg0Jhscono8iPR31pKa2aRq4d90VtogcS/s6J
PzUaqaEV9diJzpzQ3KwccW7KiNOQbM9KRNw49E1iHYLvxda0R3yuYJ11yB0f4KdSjRFFUao78Aee
4UNJu1DzbBm0dSooZsfMPOkS4EYkvY1JQKT77ps9vANQQ4UkUM9oiBWhM+pnyBcINqFqfmBQuFyu
uQWkzuAgxVa2W/dnlUnU1iFRckwVyexvMnVq1ZTXxkIfvWzTO43M385uFreRrZhJ9XKAUVYVh2F/
pVONZ/UV0x+38D0SdlQtqQ4Hz9Y+jVx6KCygTtHT3cIAbBgOk++oI8bgkCQwwiMO7qyV7JkeOlv1
d/+sp3/rJqhDeLUVYmCrF7xFuWsxlN4TZCBIeWYIfsIxD1lox9+GTSroIry4o/tboJhtieKQBxtF
EiZ5RuZvE8QRDv3NHtcob87skTt9f0kBbP/EVNuy1jcTsqmFFgXvu4t96kgRE7yep46ZSu8U05wm
jZg8TvIpXEVsnRqejRTNrPVMAm50c0c50foaJKiQNDjQQxb7d8OtUehjp4h+kGEFy+KWLvdOi/dN
zLPHJ/u/2JsvYyXJ0AHJzrhl3vYHgCXrLg4oBnuwGFHRNN5h1N3YfADuHY2/HzeCAJtHO6TnWfS6
6XBBfRt9d0cEdHausrNxE5gt4FOV7iHeXbeaNEPiMQy4DxBvJ17q8fjUq4tCpwz6Vhn9EilwHu46
CvTAAOzpQTNuJuyA4KI3kE1lfPFXIV0LszcDZyB7P0ejMJQVfsfNBnflMfZ/Ac3Tsi4650VOaMFI
ZP+0NeD8VKSIf6xwV2hcINJaa7PbvKGFfOAo9w0Gxwnl5pVQzM2CMYsJ0IJXqaI6XmfktacypzLN
NNH0MuP8ICZVR+gVEC0GHtj/OQ13xjTu+fFBimGTFYPXMvr8CQpcZbcAw5zUB5iuDTmINMBHA0rJ
XeMcHp1c3S4PlGkdmQpfJUGeJhsirCzHDLnGuzKmycJZbOyyxlDIJvH3N4EsYXYP7KsRbsstTQk+
aXpyofSTiwi5D3YjLRFyaHjihLmrU6lDxu7Xud5S2GFNwI3dgZBgcM+pZT6RagrArYVcPbRsFEll
1cstRBBMkfM4xASCvfBZzKJkI6brqDQi7zjK5SU+pZj8g5aY9U42K5B1qo2qP2fVK05KUo8c2rHZ
Nia87Xs7zXBKghGspHQPZLtDLR8W/a9cwUQFsiFoKrhE4muet4t1yTN6GTcTnIyCbfdnUjWgCLKz
UkmhB0oxkKd/vhdlO629T10+7L/q6/kp6hWcT9KDUVrTv2nI7ZIt/+tTQWA+ecpb6SBCRnNA/TkU
vHDw7k7caFMXrgkpwfcdz0xgsKtx4tRu3E66lDRmNbz/dIxzY25lMWf7qAeSb6rQHch2FxNzz98+
Aiv3giiJvdnxe3+vjzBpVWSRz9IIB8JCpI/zjWFycXiZSZfGFrznqn5v2QEJgtnlVSdyTToTjzo1
1hVNT9iiD7aBGriAiR1gUeyKFGr1ZsRu2mh+5GcYQoscQp/1w6spJaQvRYwGItkzxfushxYp8M33
LMr/v8+7xU+gF+gjkEMVC2xFdDsVbTAGwIO+gTQMKGlcqPQxOldyKBOk7i2geqkRqjCqhcDeqIyO
oLrDFh8F6mBgfhrT6F2551TkTH8K6ocfAzcTdS0uy9SArhznU4SjHas4RQquuyQ3ynoLaxgsdSv3
YPG43CPtYCTuG8tKm4iQjW0wzxdOy6rKWTjYWXciCbRrBAUCtO7KOqQncX8hNjLvgVXRorhTZILf
z7OKN27CwRX0jWMNCuOOYLGjuLitTC9G9/ZYZ3p01MazsEUTnAGx1nHkU6GnE00dHDZLg33Q4NdM
pJTQ7KjNwS1c//Ds/4DU5HxEaNL1Chr6mqexhQMACJ5fPk4wa8rLLqwXbgcYR+o6xRGg3lZARBSN
T6lSadBc1/E4cWS/aWXrxTqW2w6lweZOOhM60DjviS99jgYKHlT6YfSEIe0cSVC7dC18lV+YWs4v
Ulg/NG8vk7E8fHkobvaSkUK0+wa5q8QJLBMoxLKtpqwPiNOYfC21Q6tVRC9XvqWaSxG1+UqeXlv4
F1UZ+T69tFBCvm95BxAvU02Zb3qPPkjy6RXIlcPyFF9CsTs+EHoDg/AVqPNlCIB8Uvy5qiFyELZr
Ick/w6uEsCcLebqa3EIz8wGrOFxhy6yF0FfQVNbbQFyOeHswRukedRmtDBSndghREtivO2vbuK4t
wlpfPo4EksXnl/nziVoviE+KW9EFB8Obs3EWid/I1KaqxLPv8Lj/90nOY8YNyCJ5PwC6qHgSi+aY
JbVucpwNDo1BWM90HDvKZj0QEQ6qe+hhfPzE0XRjUiXrFElfEez0NkIVWpM+hSsQpgMc+kqfAEcK
T8YDTv9XFiVBIZVYWQIAGfoEthB/GiYOcHqjhcyHtn78LiQz1AQvJvM/L+Xgpdk10EQ3iNgZ2l8o
lknhVLIpe/ZY8UUzJuY2g+eJmW6yMzAYIsCmjz4zfpKexw2/NHvpuc9VL1en7gTjKSbf2mYJo6yv
Q4N0pPrzQuSK59WS7/jX4BwQixii4gi3t0nQLRSyvnIo8t1x+D6M1m0mIKxhE5+pOtENaC+D7i9T
nP1OBytd2z5zoGeC0k69IigkDa9YEH1oSxIH6qrCO5walwp9JrANnOHTuLvQwe0OeGkw1QUOU8ZW
wXAcd6Qz7mvbigyy8kDMW2HY641UfJ63zUCB7hit92FLvLXykDwP+uwg5xis2B1JQohEDBWzhsBL
gHkISRH/NNimsfmXUSvIQeSpMZrzyUc+vuCpijSFp0XbH+aSA0BVyGwR6XIve+X9i8CzF7B7in2j
O8Afb5pjPKbNAtmPA5ZNAXI+yrYS4wvr6BPkabLzDJlplMzIRBjdBGjgTauFExAZ46A16KSHNSUa
N3rEuxtinDVJcR6gWFITO0vPheuSZFVIbeP7hmD+c+o7QP/NZ7Dp4+Pk8+WZ3MvnQ7gLaE9Ljuov
LkY9lWxQgIX1WdBgX5VLisFhgaRrMDqV1Ma2gLZeeDggbxtHfNY6+Z6ZR/CSWuw2ykIaY0h/wUBZ
dYp3yIKAUmPur0NqNGpNd5W9ETPRfENRKNIAbXCDja2t7qL+03dMcTZHxx5HRMfVhuV6oGs+bwK2
uQbh9xHMPR8v2qxOeNxQjop1jo+04C9C+9EuA6qQZinyElOsHTWENkar+FUyAoELXoWMlemGhxC7
FLMC+ga5Oyrxkk/PKAk8/1Fi4PPRHxBA07JmIo3hLn6+e2ytFRsVFEW1h05KplngEG6nZFyDL71e
8syr/1MJNMUEiE6ste8X5HNG8p8PYWb0ew3269WSAQ1ldnVQIChbdvajKYffCEwDMAZaOPWcrxO0
Ei/qLhwkK8tzf3x6anZLXTeQB9/WMkVkxc3z/MgCvCnIrQ9PhRNabJQbZUo7ZrRERt8vV/Bkp4Vp
HQh+KObDf0acdvqrz/28K3Z7ohRn7r7Q/jhRfl2CLE5QKbuZHdkejZtU0RkbSlXcUnZqyzATMQ5m
K0iHYGmL3KuSIVtubD4f5OuWBkjTL+BAoE5wrSSt0jEgSYFIC16Cm4yeDlT+31bl3g7Otfx0tUjQ
Cbu75lXS775F+caeoYSbglCG2eF1Z0kYOg+7I78etD/rOuuf4Auft5T1OZ2znWPa9DDB9D36Lajo
x3sMs5WBttz8ZoqEIMq5WZ1KtwxSQpdZ0Je3oxz1awH3vIrRTNVYOksQBtAnoUdzbhWbuByKC1zD
jkAvUW7roS4Nw3uaf1uXZB82cghiOUPX7MpUBicJvzhjBi0FGvrpakNZfagvGMPi4tEcbmYYswgz
Vn09jGBe6kihDuWCSrfAt4kUIlQN5bqEY2MQesxN1i7uqvhnm/tQKRiFNy4FwrteEjaXDopwzcIL
l2LawQ7KKCyZmmRLgtJ6h5Gnkg1X6oZ1xrkoxWtki196UihDiv5oDNF0wRwwop1tcoKDlbpOtMGA
gR4NYySrB93AFo1+fniE6Cswtt632sxqUrY+8rPBJlHynBLCJ7lRPyUb2X3pYJRTlh7uWfA+4VqC
RbHlz1V6hbdv0eJ82DhoiQln2dEdFpvUY2P40JXAeaQmpgdKw065AjZjIVXtdy8EtbFG4zWLBpLE
xEF0lA8qVsCg02rD/+E+TH14f3O9K9pCJ3nnv0TlbVkrrXTlZZenvqm80a32xP/tVdx7uUl08+e3
7CVhBn/p6U6vNFT0U7g0Hmt7/WwaahkCu/EljKjrwQGgVqF13zQAkdkTDrORuGsov+S5HhO7+nwG
tDgJITj42ok85xCwOeHhUGRscgltnVcbFzjmRjfUsuF6ei7RA2XznOrKxnt++/j8AdpukdIyMVFr
7jEGLTdhl/i2EhPKolVlkZL5f1NVt5z4gx/jD1ovKKlDcR5opau4U6zYi8SK8N6XHmr2HQzidqSW
RXyTvfANvWyfzUKUU0gAhI92ClpHYBJcM3LZ7OLUeazABuBapaJs93UOmE94R2AhPqmP937BBTKp
mrK6+hKo9FUEV8iwPqXCKANU14rqrsbgGJrMnTeev31cZftZw1NJrO2vBdm8vuq0dkoZBOlSkau8
SXmd9E8k0lA9QGe7gaTnrZMS96P9fmKRfacDSaEpjHhEJ7eaIUKIHQ0IxBav8tmDJqVGwPhSEDcQ
SAjix1FpZ2yZwwVqRnHdTBU0eFYKsiVXrM0/Rgz/Tr1ORMcOIG8Y9mcU3IV+ysRtUG52lfVFqnEi
zw5KsvvE3LH1auagbIBcAiwOIeKVAsLPV9exv4pEOkLo4mxi5vUh2je0nzXlA7nZVZdMiHVAtpyX
KYznbzxiIYHCsUwBR5hNLJq6Zu8whOQwggZddzapqd57z1kiDvAD1iL4EbcIyyTrd6mfXTzliRYt
rwb9RJb77a4Nj7u9JGFxfpr5lZZlpVXGpjq3T11dAHt/uzIKuezfS5JlXzCnL5kzOiR1sQXlmjTK
115HNzrQFTV8ulugjh9CROcjyxSPX0rr4qtshPuxRR2NPeamwshbhPPVhxLEHDPjxjLnm5NNorpY
8kx4VHYCX/IY5AbJyftak4Xva+G21mB/7jrNftCSW/tqvbkeoBSCtzqMAwmBPAp4fuigl365bBVT
96tDXt7DKCmMu7HkiNmSU70+kTfPyjkUOSOrxwnXFP0SOvW/dvCqlE3lVN6gN2i3aEFpknQSka42
1xKDff32Sb7d/veCH8DlmH/lo3hfhJlAoVo5yTgSkxIn079+b+UaCSkdjUHlEnmk5Mtj5AAyQ57A
TQrlxdn1PKh7nUpaaDFpkcZVKmIjkwKN3BiHXqIfGycuXNRryg/B9+yMUlQQy103Kx2P24Ve70mV
56X/obByXswQ3Xvl93rCGMLV3d0Kl+paAwLrihlNmzYVEt34ANTXSlvCD+NZasPUKEPiSTEc6MCA
WpSBexN28wAPvMt7d6fvDjZvR7SXJm6TjAPd/bmgCtQMbjMUqz3i9Kb0p7VTZcDUabph/sLvtYO5
P2XvGmgVoJy77+caLK3nZSqSuPgSMGC9iut/NKvpqSJlz4MvifEHikBWPU+m5Qm+zL51pLkqzr7d
sULR/PNGyqiodqzpJEZN0+qqDd5TNT+07W8QO5B7A+pVf27XwRvWcF9thssQoxpbReUBwt0A4OfD
iSTNtwANaZqhFmqxHwjj8PNJXKMAO67hSauFscpA7VJjYAn3hoztGdP/uSrl8Z7pZOPujidRIk86
AXJwglBparjnWIwqpsxsQcTZVMRpwyqFJZg9XTuHlmgSiHyVvBLOAA9ULghRa1XSYJFFsR2+APpR
85a2D5hnOYsxP7dE6xOPJbEUm0YoZ/WKeuUW/+a0RMOTNDyT3aDZ5YgLtYT3snNtRl5ZKCWa6sAC
8C4gc79QB7+FljB6LBRBbpB5pF0H2kO/jPMBDsxEMO5ZS1byGFFf/3m3EHHbPSnr/bLfOTBm6W4R
t3DNa06tpSFJWKTlFLY1TvmpAc/9ad2Mo49KNfmyVpZ+tmtYPok6R5yy3JW8mwg+cTTeqmWfKYpX
V5XSBoe8SKMuy0XIFTORHwP3eBTywpl6x+6XFMu069XnkDXBSuQCXqLaiVIwl4wDjt6N0DLA5Wvz
RjMar3AR3lpv0mTB86mYWmu2EAPMrCcsvuWm8Ht//9E3cgkuVA8Ba00HfvXABJbr2owGStY7QATY
bVHz0xicAaUW7vH9Bnz0RQBdroP4eLUyjUXkTFKPTbuveogivifTnLXM5fuoIaa2rAPCgf++yzPU
yxa/cxETfyqpzYg7FWNFUcPF2xx/S8WcpS8LGY4I3kYk6VJQvN8OcMxnOa3Wh49f4Izo2+HmBXNU
8wwp2gtljKFl7KhEowBgvuN5YAKaPb2aEgD/KBZ+Zuh9C0d+EokREB2pNF0JnwKb6uNHAJM//muy
vgSGvAL09Q7LasQ8/epxs3XqDFamTpvYKBM/ZghXpNVUrDIppExkx0t6gEWf6DD89yAPcIbbjAQ1
PhxYJeRV4Y8wz1Mmg44W7mEs7CK21UrIibpTlwn1+vBBeAYFNHCekRMqkY1QnEEPyT77hMZZ56p/
vyq3ItvORHNaS8sSvyy96xYPiIaHqrbPhUQPbFJlbL3EnWsU464CcJ6igBwFGf1XgRJ0F13haQGu
4LaFGgJ8NH6SrECqZ8BGZtZ5CiGs0pw0BTPD4hOg5/pBL6yC33UENvHFZ91bPTAWnmaJxUs5hkQN
lFZf561zep/k6EtPEYdMY8MucyBjbZoUxWsanzdYwgJvtu49+SHaOquRBXnaHe6Fpy2sbp7onIhi
kai9x/f6cOZedCiSoEasyIpMtWtUUwqBX4sLSfuw5HGC5vPh70frNYmYsn5E5oeDDI+JBXoNs7cH
qyf8SxMtiOvcPz085/448qsT4j6zYpmeLXE8nr3V49eEICEBjccOi0qcYfEQB0AKqMqqKe6rCvaw
keAsdgyOc65fA9VEk8aQCWiNrdZtCp2ggBrHP1i66rWwISE1aNa8ndqpBXBz2yU0bhAlvoLyxprH
uzD6GMXouaR1eJDjJWA5SqWUA8nROuWqL9dpZqMpbfzqAbHDGHR2I9wLJGEzX6w5SogkSekcirIC
n2sGRl1jQJLD1EuzcEYLCRBrOJmE3LKNVPuN81czhC54UD61a5t64ba3kS+MLm1TpiUQ1LqE8oTS
vDNAHBo5qwEizZCMoi3qG043CCO52XEuBY3samOrMGQEA+47xGezJk6QrpY4ls5u6UaqCehQxio7
W1l5cq/8xRGd9HpwqRk8Eppy9qxGRgMBdBEIdCAufrADBepqjh8pcOXH5neAR3MrQXDdn77fM7Vc
4xFt7X+3VEL3wjp5gzjU+w6JRXF/V+/XWs01rVhWLU2B4YpYTJTL+q9MmtcUdpvtrAnr/Eih2ELQ
3XKGs+cVWyt15C3tUG31l/LFQuqn+xn7UCntTJYcaWbhBzv6AAOui+9xfrBU9/aZf1OORJiuMh/f
th90botj4wqn2TKZbpgje1CeR4AoXT2EHGnCrR/3C59Cc/Gn1OcVCExjBqJ43Dtme70ENWK2NlYx
eyIaUeh7Og9XdJN5jkKmYj2Y8vhQWN4nXljyzmviA4mTkxIEsSPL1AMFRKPywGcH+7X3O+HO//bR
fg7IzmOGEIJy2mtO+BphJ0Wo+iV1efuLrfM37iwqVlyHLpE8XF8/lSmUXT91f6wkj3xNy6Nmp3fu
oBpI/PE/2/ypP1DKfgoIyhgdDvGLyeu2yKAKA38rWdknXyW8TrL+INLz0w8fNf5YjsgspwMjS2ym
z9MqqAjO7ulBAt//XGR/a6yE9DzheLjzqEm9cfpKB6MI7nOgvCCve8HoXKegrlW873Ob4nFrXmz6
SZmSyTVGsAX5q5qZvaomKmmRSoB7AAwbXwCyacEHcloI6ZIBQtwzIKuQP9Qs0tOaKad5ypPhTjoi
pQ2/yGHYY7UtgEHLbGQqYJlWyN/6aime8YNbk8GnnwRONSGflnrQgrV7lj2gQjvmKusdJg1nP0pv
PzZu4Um5R575EY2s+m2Tb+2F6ZFV0R7h9yZhtYZHb0L9kEW2OXmr+nMKvu4IXiD6IVSLQY6GCbfY
JMK3OlOOQu2CIJ0cJSQGa1oRfoCoKftNztYV0Zkg5CCROPk/EDDMnzeng/r2DsAAyq0NcFWSFAuo
YNatDxUETqCp6MFpGXGK1pngUn//OAz6ncLMD11272REPf/g+5wDJNncc0iDPQd3V7rxmunzQ43a
LHjZGlFVfbhKZaE3h+OeE0FEagprgKOW7wizxUmGjyQSX28LoIUA75gzbu8p+pd3PbYDvVIC6i+/
8W3JBTyBqEuMh3C317KpYXSIsWUbhuFdT7dQd2KXJoKGmluNE0f7lRq+bRH2Fgy73tLlxMWPREZE
cA61wlrw/oAqPJmajKlcQTDhUmR6Tsnc0QRb86vwyAs5T6gt70eIYMQvXp2RRKhzkwI+fbSO1XT7
Y/Hh8JlsRBk+vI08B7KMaCTirBjsQAeL4apDumuyg61JoTYzFMKVn4YN5sNu/7KuLPpL1jYbUNlY
O3L5NCz9Cs25OD/bTlzO4vrvyOMIXLguI4eIg0b/OUE5JbCwteYmitRBA3lUtFBZ5034/9dNuHiS
+01lCHHZg7O+bDvr7QYRbf7eD6uvcOAWug2lz38w/UE4idK30wMRhr7clmaBOgm6JKOkqplGFK1R
C+XhMCC0oAtlLXZcLpln9gHxi1x1XO5MNkIJNn3QMAA1p1vdvm1fzL7VjiWzAi90NAp0s8+7mhyp
IdpRp8pPJ+E5qsFXOEzUsoqOgOpJbHK/QqEqgUeh6kp+MjLiAwQXELWROqO2g5EVaDiWTHJZ2mfl
TIgJM1vWu283uZfjYGeop1nKO07lHbWjFJ+eXVi9f3QIbfS89/Ic+0k2xXkcgjok8PRuoOmlBl2v
u3oJVvJN+HG86AbBbAUbahstKYgndksPkj6uZ+WwHP2vvGF77ZyamWnT28ZA/LUbi59Yl11juKof
pbhRjatKSTEnfqO3PBEisvc5YoV4SxX1nEzNez8KhkXxS/YKQYq4/vqT26ZQ0FUcBQL7DwD0Tl5b
lWaY328xx2GEfG0lfzB4wYXe3pWPi6yquFJsQIX1lqPb4hz6jPYjbvilN+DaGRhjpYMXQ4l/vveD
EhfBbL/Cm8hoWUbc1tsUDEoIia5g0pwDKmkrUTC/wawoLcQVr//AOTUWJj+UT2nF3ZAAABip3Rap
Cdi4TNmLKcbnm/yCgDfQG1uSF23pKsh9OT4wfUbTkdbfvSevrpL3ijajxHGxrhQbCRHGEUFtrcah
Dka1TpqKOW3DujLgxV7fAfahS/aNRCYud+0hKD/s595dWGj7vZ3ftgmnzZ5TC0Sa+QohawrUnTlJ
kJK6QPhnLC8Dpl2V6b7fjIdS23EudyNIM0lEMVfG0jt29jSm9rolN++2Dup0yH5bxF02d7cyheOg
oPpSZSRzF66QSQdzfXJabFVJVB/RlV5Vrp5B9dj+LrFHOaZO7tLlL7e/mPMtTCYPAqLp2kthYCcC
gD6QME0GKMgt4A8ukOhCuZj1bx/al1TNWfyWSeLamLOTWuvbkMQc9+aD5uX41JXVgEy9pBVnOVg8
gwKVnXFb1tq34CY91i+0i2CPZdeH7LpqINX3lBqbKT+ggZzP5cj94fIlUc1NUbXQEJY9E3QXhl79
3TF/D4pQZAe6sXCE0me2M8dWrVdhqFfeKiyb4UISpvCL2KJ56k+eviU0W08okM7+TrFJ+tqNtiLQ
IwPbGSkigcsG9b9wktUacRjY1T65Y5YIhtOWfyhk38WxXJUYwG2+qpapxzFCKl40l6s674yqLzVX
v9pJMQskH2Qpk65cPItMmTJc0NLaIQFUso6idqMn4OEXAgjd+alSaMCWl7Z2fbCU7ThjUCJL7xeE
XkWANBm69QF6d3C+L6Lp+Qw8mht0ixs7n0VPuTXUFtrM1QawI2Ok/yzkdnBM1rEZBJAIRZeFiZOw
/WZuZlTIvVX4uUuFiD5XvEb8Uyoc3VMiwT5aSH56dPqXqap10RmkrGRh5uFbt3QkgR+Ja9Rk1Vpc
K3zf0kM/4/kNODX3Q4VQIUBP+/BMP74i7SahLWE1blzp5fFVtt+HK8Jx//Joiq0QkimrM4JbnskO
8NnNfAG5Sr+WGUHk6R/4AyiPpP8Z9Y9R4Mocc8v9JWalINQixuTa0RvHHvyWZ8DnTHO7PtAFVmN0
e10U2fMGLozA09S3Fi0A8RfoQXBX9C4DxJxj+SZ3eqX7RWkrwg8r79Gd3ofX07wLpQos3vHi8mpj
UypBT+REmPNYxXXvwwoHvcmvErYCvRMem1Z54LY7t55JqjIkedioP/ivnLNGwVIfLQB1UnwjWF2f
b6mtCwjR4MonxORqWpa8RgtQnc7ehE/YDsCtJ6lEoaksX0kfMbtevR3Ca3WKcvuIjbqDSU7xFSZy
O0GhJHFrsCWEtSOFQnwaINCUCraBmek7JlMX60ZeOQy6wZ+iZftKRC7XhDVyDvnt5/dxyhTiMzev
7tjz1BNbf5D/XObTie5LiKnWdWypiIDX5BcwgND0wT8D6C3fzEVtFaTaqxsp80gXlg+3NuYPzAgn
IMY2p1jRxW/3N6by7Xrp1RtqAO2olvD2UZZJqlOknXsNN7OyuM/bPVvnpbcEHiOoSaUt5M4U77xy
uKZ0lwlGlEjI93LjCZm0G3HK7kvtq8DFsI0EG+/zLJXjRmRir7iDIy6AhT9hLbzjZk9IfZKSTHRu
6ZFczpMnpCu+aEL2gLojRv7ZattoVyqtljR+kLRGTRPoIh08uGb/AAJPtIqfMZGh6EHoqqTWcWp3
dcj/jIQlTVL79o5v/0aMv4McM0kD/ZPArPD2onSdAbzwuFuTPA3HaVnMZblQ7aEWV+6hsET9nq1l
S0r4drz8e834VVheWHjmar77pRcin6TFyuBW8jquvSEdMlDCJyG4dEMCc3hwSG8IgJVLjG83Hm+d
z0AdunA6CBxqKZyddJESVYjkzDekQrflpb7pcKZV3LGSGMZk0XF2xwdVilro0PsRFoNMvhJRCNaG
1rNAy49Mi5/b94ivoIQzmwxHQENqYda5uIfyI34CeWpb/GVtX+2MbBE/V07AQWccafZvWlo+Nm7G
fCIacfg9Zil6ZyWirX3KTe6idzaglKtXrlXI7aJ4GdoPKDmtX4hc3ztQWM56BO/ubYSrZIEGO46z
t6MiPJ5eT7uCf2ZOE+Ng8sultrzl2ikjYTjbzQzxOZw9j36aRX3hi+uzGUkFAGw13co+exvX2WQF
7w5iNpPJgUZWVhVbo49TIpZYKCX6QUOclA+Vv+LmeSIbMT1djXZT9bo++8TZQk9SDDXTwc3V0Z26
RimW59/ixqKhwGV6NykNZCi4MmLYnLjEz6ef8RgCi1+m68KSqp+f/Wx9+vyxCrb1hLJ4E8pZqw2S
9y5lkKSo4eSwGpD7N/vv8Qt+tLgUPjclG59JNrPOTLru/utcrUitzeDtFVwAXEsTX+HzjsmPBDot
o+1pJOBDRc/iFG52gL4S8ZIfEuWy8EvSXAQ4HfuWrxug0LQ9zKhp9uWNYJSCoConPUIZHK7axLrP
qCoMOMKd02YLC3WtJs+186/QsEnAfQM+IrFYdLDAEs5l++3Gusg+JFO798hNAJL8kVkFoOntR3W9
T+tBl0Eh61HKKeUFaoNxYDkZ/j4KKEkcKitKbDMzMUMWaGLwMVKOPvjrr4JAautxiUoGligr2reP
5GVE7gmOmc1WscUGFHBh5C9v+QvJy9lnqEb4TLgsu+5wwgAO0jjcKuN9UN9iLAXEYohJ2w3dmTHN
ShJJ7zM3gbRwhuBdDmLm08DexYIOruYU8IIfyJmUu+HWV8LfKZwSKqrXkl0kXlSu0bduLC8JFH/b
dmLNBv39OZj8bAoTu86Lsa++tGh3YJ43h7RNdD5o7HP25gsUc81d8HGv+Q9C5su/D2/EmuFCIU9Y
Z7hXARWbayeNZd0kgctBj0ZRxFtoiWX5ve7EbgLvXF1qdGOL6l38GW4U5orAshbFGOmG8XQ0TV7C
kFdjJHouhsOhaymAG02/FI5bnPemDtAxKsBB8qUmT731bgjGVYTG3IsKJxRdRCYe2BU0zu/6nnM5
axHo7SeW3FHsB5oEpkEmn4DkNuaLk3DU+IWl/znymuzwxW3AMn9A8LGOG5m5da6AmZmT63osBqcd
VmRtZon3KiTPTmXdIHu2wWRtShAAhZJHplOBjTfqaJk/FN3bxqiv2ooTeUGTGRJhaab5J3pnJRpY
SgH7NftOm9Wbo0WP1JjjSQYq1W4Q7h9cxOVEVlaVmCpFt6QdTMod1+5daR6v4K3LcylG9PkE8mHw
PgF8oCm/q2pe8Zv2PP9/WBzW5FBgNKLcHx4P16py0XsH3k9zDF501tITEogWwW7919fuB4+k6IJf
WKnPKouU57ojJwLcnCTaqA/FhiMW1X5v/6ZWXf13AKutFrrSpY1DI4eP7Z0d3hT7+Rmpwwr/siiE
FfN6E/CLaI0opC0piHKOir5ATEWNgfdWs9V++HSufrtQQj7q6pa25RQFoa37mesOCik1s3bmVAH8
sSC4OJT5CYaOnRA37G/bgbzbMMykY3nEMwCTQvMdxAxtzE8VTJZoXPsdVUJdLp3Z4kDuGkGbtcx+
v1ibpxCLMXMvegMK7Q62u2SDLsje9IZ+je/JB4kcNI+i3+BbW9NHVZbr4Uk/1bLSlmQupzt40P75
AwKsybfvX/qdQlCrZHmJP5m87XRnRkFXhajgpSYvrIvlZkmLksZUMs8LxoamgwptIjpiHaFR3p3h
qAqNCP531vw2vPsV7rkEC+xigAofPMLhzAKoGuC7m1DDVG577/iZFhJcgewONrUIbMQ8uUG4o015
7zDt9ysEQXVfTYDzXy1NR+EyhC5YB2jdFxOSSFt4xfEAHauGaSpf/P2FZe0zKaKdVDfDvxymfHpS
VB/xINxgHlnaOZOp22PHO3vCmaAWyB05L9isifxD9+nCVg5hYf08oGRpLK/Lvvd1DXOc5BdaHAd1
G6aA2SuEOBQeFzu5Ed9LunhuglHtGwAvNl2hIijRswE9qkd5kV7m6e0zGjxrmyUOY3FXnV/bd5MI
1IXaWMT3pRszWD7QqiwpA+GvY1jftySaaBkJcUDFZtmTDbE7Nl6xO1XqBgiU7+YGApEUngoQnBL5
AeEFUiAMOxgAJxqc6WZU6+UMBpsmEX5neeNlOdzCTCyeWipf3a8cap+/kTZdNtKvRpgPTAqW9hPa
Hep0nBrpUj2AyhYQZDdfKnZhA6pfTaLzrvKq7W+edT0A82KdaneOfmGepq071CtSBOdHpN5A/lBE
5UhtS6Kg2A0LP3+0dfT03E5Aai++8pCBUqByAjt4lcmZAVDhvFftT80WPRypeiKXaURs2YS662p9
s6jW5ql/ZDTw+OfAlLk6/FrpxAaUxK+s46o/Nt0EH/w7KJp4Pc5VFl/Yj7Lsets3eRPp0y7GRyWT
ecjh40x4d2+I+ApHtjfA09Zocv5dqKGLm1e1CpRQShDB7NQqgc+VnB7Udu88txxeHVuZ8+9paMXj
Tw/hLnfwUe9kgAV79dGS1RH2/43G8X6O00lNy9CbBiBY42s76LuIcI1PWSzCI8P0tZ81/1uDcXd+
I9Gnm8iBdx41KPuH1HPG1A7JIMafs5f8Uq7quo04C1AYeBL/jLn2oCZz/g4lX8IyQKkeW4kDO75f
N7DBKi7uDt4yCJWMgJSauMbhFYH/k3XaHb21fEx6shYqj4knAHo1HEeBvmlDYRuQ5VzgKLI41Eop
n5bpDCDS4YCwlGrJb/kJ9iOeF6jbzBi8Kdhk0Iyfw1FzsLbsv8nWMzkM8XxEBxZszQCBZsXlQOcC
CpiZXtMgALKBMv6aineGxREMX/1B9X/vHtEVIzRG5lCZ8DO+vRcC3SE+49w33UAi63Yf3Sg/idrg
hh/5sXToxQkDPbebpsg7PJsZvZBwQgJ1M9A/DlTr+Ww/hn1zXHgFdz6Rpt55kk/MedL963KEzcuD
pYsyRRUJjjIT7iMCvi0SnYVESXgnVq1mMzckFe/G3n3+OTMbIe/srsLnPQwaCWjzOZkssc1iN6S+
9Ec+1c7lFrokdRmFbZDiodFtES9JbvQ+HoyV26kBTtbDG8pbVwwzKUW84BcJoA2M4Ou1rE8Am8jc
x29/kUWmks2TDIUrNvz8956+Fel9LVGiSlExj7ZwX0ho9jztW5TG5enmE47Yqe2As5r6STCfGU8S
f+HnG2/QEWLHcuzEpjgoEDscArmhFO6i38JMXpXyM4/hlyquoUf1pMBt2AkicPZ7hd8sr3d6hdBI
4um//v8PA0jLX/kZ7Cmg6zp2LkhRI9Lpos8mMg71LqjOJFIU1uzsXSeNBCRaO+RtBzMpo02a/UHV
F/jBCyjmUfqK2U9YgDThlxYQL/Pso3tuQEZ/8mCefB37WKd9UZ5SQtf/ie5ySZPmb1QovuHsOQFf
dOd05dFUCyc7046f32LbfuI1Cs1p1jYzIMf5prMJLeyGUk3fnsEtRIg7iDAH875xt/BncXUAjrtb
M/cwLne/0/a/IPWg+ZrPa9Ky39Oj8IHd/HgHoHayHyJToRNJTuOkBjAcg5OaW4rGqwyPs/mEs9lg
sA3xASBeECndH06R1XFB5G5Wz61q8FIzdTAMUmHnvteOm66LyLtgwv2yDg0IRtm5R/RT0UxM3Ay5
EKLolApeThjEVjz4cHASZJULjWU/XE7uOYdfspu0Asc7kKRDNXXJlAAN1EbWNTyXwiaVzjpgFsmi
0k6thc3O7S/pa5SkpnGLawidx7VE4ABKi86hAcS2zXzyH0SPec43X1jiCQOCOByH10EmzntnB3We
G0SJ3d0dSnPpYeMuCYCkPJIkh8NJM7fYKu1j1p2zzEW/7pmP1xXLneFHDK19UkvzZ5fZ8VjyeRHr
5p9yP+zytJr517upylX5fKNVo+hYWRx2R6F2OdjrozpLyA2dfomumZMh0Wvv98BZuY23yw8LaFs4
2h1MKmSce2veFhPaxepGKKkDcXSE+dOARd+nvefBQSZ/BBnvGcYqIUMr7wH7i5kpM9FVgKNSCRG9
1PFMutceov3sTqbjk9IONiEZLu1tnruuQ/KxVebTa+lKOeKWIP2Hvd4KIDqi3UauT+Iv6dNNu92t
/DwDJpN4oeW9yfNCrGoGUgvwV08j3VeY4WsSv0wwNgYrhusTTYFfi/TYP+vb5IfzSz8G3/2ojwji
xHasJc7nLTMWhWjVurwb8+1yJHWx+wMx8c2OTcwMm+vj/DRM7M/0kLHwHOdmSKCRn9MgZ1vGx6Gy
KzR9bXo0PB2Ffv2sd1OLJr+IwwrrtVg8+BSCE07z3SLZfODlXeXG5fihSak3t2aeubn8mbw9stVK
nscUUHlhq4zElm4LofVwsxsi83bbZtkUOpvuUCxOxSaMSypwpARePG5mQm2abmu9e/CyA/jc+mqO
TNIU6pxc06GbIDKZV0dEVBmOb9IM0ngY/lR+MKLxQV/3hMmm+vRF4xKb3dYtMZLphz3fxempu6Ry
0z+cnLg4aM3+4Dy4eA1dZihtfsSpv3eJyjN8b2a+HO60t6pXaf78hgtn9nCB1Tb7skN1vzSEEt5H
sShZVoiaXm+dbKg+PqGshtdJwUzLk3vB4dQYftuMOBPkgl1HwRqhiemCpc6sNANI89B0zhxm7Dqw
pxY4En2USCWOoqAqLZ9XHoEjc3PpfXCOgepBJs7Rw/ub8z2JYLkxRTO5RTacxXHiyKrWUSA9YMFn
DcBoqIbN36wn4l8MykTseCgY8XiemabMbb8VgxUscJtO8by/VRodCnCRYvvcp6A9IbLR7p/JKVUp
3eJeKVagPtqZ+tW5ZHvlHPqM9p8kSrLoBQnFdrZDx8VeoHbKLkVc/+nlvSxUMUEwKF+QyTDY1NhN
OY4l1pCDIfaTetrKNP8bW12SP/6nhDUfS49+2sm/r4MNfoNJjCxGBiDCD5ybAFJ2MwPr2h9Ba3k9
V7p6NIoTznx4LTt/IhZqSy83gQU9mFuBqiJqRgQ5z1Ck5mk7+CLUSoPNJVNDWF3QWR5WEKFBAZCq
9Ca2cVFCqH8y3NM8CMS64y8WVyJHj04v8Sazm+ejxf63IrH98d9eutpT0JsTCQ3j5PORLcMawKIW
vR9STOuJszmjDr1Au/9yOangKbj4HbAwo2mxFPIU4Jdx94UREKnCYeEVSBkNqqMlZ5ZkneZkzfMx
Q41dOA2jiTO8R6ILgZitWjySCfKGcrcUFzOZ/EVY3E2FM+5BUWmGNnzCe+F2ZXeJhKlfGaY+QzBM
724MGkbFaLGor4N3O4c9GMsD3ES5NeDbu8DfInT5pLl2nLciD+h5FaqWVGGsfBrSDKum+Ii/oqrV
k1wWEsiOCNHF0jjV8hOa+KusHscB1U3v1eDQqtzmzcx9BsH7vW8m+fLiYUScSZTuPzkGFMVXViLp
G7+eYlzDp+ErP1d1f4IPU7Bz/Q+PJ0wXV3R7xJd1ZDMArBGILI4gDnQgadUGE6uMFmTlBbiJe0ZC
coOpkABYNmlQihv+HOs/E5gvmyc3OV8emIv+zOJc+a66PNFLEGYPHZ/4noOzNG1hg2rza0hyZYyr
VZu8iY9ANfsLHJTNAOrEyA0WsJLNfAXs/XybJnYKsd403aWd+duu+VvI1ySobm+XUgTI+Vg4Mpxc
zOlW9cLgnVOwUU+szVUgs1IZNjnrcLn3wKXyrQt7MHgUPcs3Si2hWfbTS1ozvvCN9pzCcuQlHwvY
GjRbOQLfIsOLpZ8LEStZkO3XqnRv+GU4pFL8Fg315pdxDr8K1Ex/yUWApwAgsnNa4u2NHad6m7Ql
8VbQLt+vITTneQU+3lNZM4Z5zFkxtMcy0C8zWX8XQKLopumUEWIo+HYtIcKxlTqmIfMeuHEKcPKG
256gZvxDGn8Bfzh2iiw1x7OsrFnftr8HNwxTZZQQbDU+PfmGmwHkWmfvUASItQx/WmEwH7xBkH1H
FSjlxbQwqmkkIZ/7eleaN0CkT0BI0gVuiqJg7jsQwi1UJ4lNBp7Dizp5sWoaa9XJHx1WqEn7qQkC
S/U5ikJBPckJQCUo1jYxgy/PPpgMGtxCqrN3tzhcj7PVj6az8qICmabpMKCRi5UvRm5+mpNIMnqP
GuB2388aFUm8wFrdPSCJSlc/GcHtj9W6Z4OQzRm9Y3wd6xq9YCBQTPuCG7c3pCjeanKF3RA38gwZ
h56o9KZq7EEKZS3LS2jipEQJNvMerY/d6rCTRQ42kE4Ho/3caA31SPDGXSYV2DB4D/nylr1p1yL0
lz2ZmkOvaiVs8DlfyZKJqsaY3SJVtWAzmKOntst7YymmJdEgW4yMrzkaRpWRp4z9V36tj7eIXfHV
aOuprX91doeQnAxnxvZM3NnmHaGwvkz5lEAqfCzBzjZb1jzTo2GK4MyLNLPIymGzq0/Qw7XQ2e9y
84V7x+gIXvgwr2ZKrq5QXM0xSpSdp2WhqlEhisxfaZwF4HM+lQG05hiwpF5TnOnbhsVIEKT07oK9
Px6lD78WYfYtqBhLBwTuHQRRkx1A0dQu2YS8YOFJJRNsxSGcrl/Ek7+rtkOLPzO4XWWkzPSwetfM
pHzQ+geqcx97tt5kl1WlE7Na/3xrYMzyr1JPH+qtzcKAC5N+FZa1Gce0XUR9G0IH5mI4WBvm6m+v
QGas6f7rwLCGpxUVmb8mc2vw8w9lB2Kl44lOOYhQf2fZ8ykJj8GTE8Kkmc81GiNYLsTsKMCBYz5n
pR/vRMUJ8M1cYMavG9BaG1ekqlwTMfRHLPpI/IuPKfwQx29OaIpd13Yhfoe1kjBxLuec/+u3kesM
HuJJApLrFWs93n0nmwhfZda0pd/WXgHWbvdr70sznQiFsVbRDw/bpbzm8Gubp4nxsyiZ/0pjaDGh
pVpqstTsZkv6SebezXCP+qN1nu2Te2NuNWSBud+KgYfcdtDj6zqdv6GO14ItEzbU8L9KGHOvqJ57
LALvb1n3fmeTss+EOZ9Etn6Emho4CTAvO0cddCnQ+8Ji0u5QZ1cwVsfmqCLDorm1I5yr0aTgej78
CpmI2iPQjIvriL1Iv9n6wH9FzXw9381LmZAj2Qa3ye2+DOnWcIF3v1UwpS2w85a2Hzc0QCHYbtAJ
jNfqk8xDzIeVPHW3cceFDfzx6PpEpnlaGtReUmHSPaFO6e1SGq3w/LuQgnUdAcEp5wbYbuNXMiRV
V4APcuoRtuaqUuEgPVVikrFy6cu4Pl+nBx/3LAd0Yjs8RkCv32gW4bKDvAerDg46yeAb7KUI56sC
hSoHOzjKwqS8Kdg1EMFBk9mG9ep+elu1wWncvZZZFHGud/QXO+krWGj+yigss1yV+UJHWNpSL3E+
69GaXEnkrrYKwJP4ondQdMaYxG+zqCLouPzn57le6d5lQzn/YtX7WnvmiwdKYV3hrnQVJYTTBzvE
IFaPtp1Hgv/MIecTmw2U8asvvdHVRJLICAGDuxttvb/eERPznkQW4DMOYuJ8VqIH3eKgRJ8vCPAL
0Cz7txmVx78n1iCRfweLkQD2InufGEJYPwhDdmfOBt2sgk6wjU33AgcbrnR/VV5geuh8NV3PZV9S
4YtIafxXap7pU5BMzjfVApGd1dNxC9r/ARTeCGesQVOY5roycZl/UMacDgeKMN5nArkyFEO852lt
2ek2ScMlTJuOC/64Q0gQgEfT/WIg0wvIA6GcwUcW1VJRpLac6fOgCNdBA/TVJNan67870Y7j1k3M
zDDvWsGQ9KBSTYeXDSpNmkfYJQ1qWjyQ6cdm4fluCBkIGskDqAy1KYY8q7V7Zm+twn6P59o+uIPy
K/qCPtoPk3pcgMXvmNdVU112hjBBFSmPUG8/WZnDFokjNLFWWPZ/X/EWRQ95hcAEyKkYJEj9vFYC
lYTgAQ5P7nO+U7TPtyKPT+CP5WEHP0t7lTgwmG1LQRREZO3U/klLdwTpkfMogsF1174iY70nL5iq
UNAl7DWUM7ROJTj4qNFp81fS/jLy4PQz38OAAq4vDNbocCAnXJ+iRZC13eb+dlhSWcu3wtmXLiFS
4VkXKRXDMExgpaHEOwlNMavxlMRISd1Lo02/MGETARz3mHJ6n3IjMiXplIzfH7KyXQZaUU7Vh2Xw
/Gxo3ZIn3VzmKJ///dFIwlFLzQNqhLO23A0CH7gPFWpZOXxxHARCPsmRvu58R/TfFCGClXJZSiG/
qcWsr2rB5AESXi1wTjJgefRrzNaFwu1ZxJMVEs2f4DdxfKmez7lbHSuVaucRFLcGicHJcFWzrnDC
wwD/KCPWy6ktFokIRQJmvf2VQds9+JnHH8CyzX7JYYy5Er55V4GXCpW4/NbeujjvG7zZ9DGW2H0u
PEaIi3o0ljMjZpAM7yVvTpXzeVHSoJSexq/mBHW5eR0cHGPqBfnKBhXyqOry5RYn61cnxFXjy1Ld
gmm6TV/XsshZYKxF3l4AzT9jVpMH2Y1t4jqxRMSGS6XaOV+Z2xbFpnxd9OqgU1GcUBigWkr8C52S
OaMbM2otKG4oWGqrc8JyeJRYqhUk2r+T8o2AZtYfg2wH+MOnQK0J+o9JT7iRLtzqDNi6Kan/ynkG
kZm9AKvOWV+s12M8xTH6oYn4/lA0bIrPKGM1c5FiryAz0JICddzoA+GpTD88NZhesbsdMae4DiIB
i2bCqHpm/YSCf28Bsk/63McNTGZWXFvlEYNRIPbFaFS9yICQ6buz9Qdismz1mjZlNviaz2B19RFE
R4eDK3iB/mxu2yCGpk4XgoeXv5dDBM6fDYcBnVzYB9nOhNTO/ihAZQ4CdkCUcZHI6ohJZaxVuMzF
4Ogp/kw8GSRW1c8FE6vaKTHL/RX3ifrn5r3hxZ8DLpllc6exQMj1G3DLflAjapoQEltqRhpUP6dl
t1SzhRowr0fDZkCQZ97ySpTr2R/9G4gHKrd+b4OhQ7POFML423ZBlbpSmPHYcWgjQWCSnHHHLDRX
BPIVKmN8Um0md7rtQu5LqYzO203nPKn1+NVMXHqF+LT7QiJ3AnAwtZ0ofY08Fq8Vi2rE1W0sx9Xe
m5qQkKXCdmcvu0Zc/CI5WLNpccKxk/hxRwbIiaROV6mv3IeSqfH5GMSn27xhLqGdQbD7Jwd8rgrC
74u7xLiHs6P2itmDj9LjYjPdK7dNA8HSfoWZslZOjqIGgugVfXyxf7DDLj/eVCM8/+oRmYoktOQd
63IvAbuB63zMazqo4HTSxZNOcovp8a1muQdYvENmwL5pD4qiMvhBqxsyRy/NQRYFB9fvADBF/neL
pC0bPdf7lnEer93PR658eqchJK9W4c8spihSnRxQUcemL/N2hvxYyNY5LOHycBIII4VCm4UP9JpV
OdW5goSc6H3cvOnc2rOOUuFzRFdTNwDVPsT6cDGMRPmC/lSY3pP6/0/2GCfRi3AAyyFU5St28dU7
Wxr8sKw/YBNDvHhbrH78mT71jk5BqSA0gh1dXNxxS4ssXrI1H/nOI81yfOgHu+0TpyFlkYO+dB1/
efpk/e+pZzuiFtGSVD9bUGCi7ZxDVX4pSmz0c2v1IJ7dA4J6Yr6SohrM0FpC+7dGHSB1liQ/KEaF
wDqTbVJHUXVaKG9LI7USJlECqtgLIqY2Bb8ZIUS1zoY6j7UX6U0q+66qCInUlDd2VfxLDozNU0/I
+VzvCWdn0cueh6o6qelIygYKPTIUEzTPJKQgbwwphli8LHWgW8ZfbKEJ1Hrw1tzZqe8U8w64CLkp
AKQ1ey7aLUd8Xtaog4aGGojS1/ac0C5djLcVW34l/P8T8ZjjNkL5eLXnsj28/L73ueUAtHuVW3S0
2Pc0TtDqCBHL89HIJEJWwLaEHq2SwMWrGNdAZeg71Yz/rAfNzo6NplqEahhhyudPdVrQsDWSU1CR
54iFKD3aXcCNUdVKxkycdQ+OeMNgMrOt4e68uyj6841SMvbDYj3mgHFvPle6mtSwyedh8xBJ/Zb7
ThvUQJ+z29za4bT9/bT/a2szJdWwZn+F0R0MUd8C8OpKz4F0tLsFeYJeCP/3UYAABS++MzrBIkEm
Q9M75/8bopzlT+Fpm/QUjKPPDuCIeXLtlDJbJJUpCA8juWHoyoeXm49TFJHr4jfAdM9tHB570avM
suI9u5GH1L4xaCA4NEEvClKJUgy7VeCJSWNYK7A/oVPGuq+vbPKkhJWsSWVFLkOIMUaACDG8X/cQ
/+qDUxdOfA35Rt/m0lTHbpWrLn7YuDYlhHswfqkYAjWlK4AwPCRyz7VSB3wzjsyuLcqLhyddrKAG
yXHvoxwqDc3Komrb525BIuxB1uGWXZ+Cve+6djf8iRwAChGl5YXZ2WEPoUsFIPkW8bhK3QwCsqt1
SuTIEHR6P2CNRWSBhmU+e+ZNbL9wZ04ZOMEcsIscfP7xGEZcQN8MOrf9c2getAUNz97OtEBAakOy
JmL9/neMc/eK3zNXo9XY56R/kI/gAu/o17iafNAfZ9tE3IFB1VEJQKh5iO5hTXQwgBSwN3KCHwEu
a/b46SF1fenBYJ3s//tS9yzkuEYyqcbtYzeXHr6AQbKzD3BQwVOIEJjhrkBcHJkHXcDevuNHoFZA
lRrLc/NeUcf/As/ygYpIVYrHvcpEKO3LuanN3xKSrDDTNm5J/16+b1PDKs7u2IYwzwmiaspkr8NM
aTWC0W+n0y9zesZ1rL1AlRrJ+XbKkX7wLvmyfgxRGjm1gFGmoEd7MMi/qRTPtLAxWzR++Dut5CCT
d8HsxNYlPz+J5ychSx+wOXq/653u/h4g7h8kb0MUFIDUQ0ZbISzyR/FdmYpiWgLHtaaOFZND+vtk
rOcUjGaEJCev42cF7Ha7pZLFKJyqp6AcNPToisTMqaacyLxrxYsMASyvMTBX1n8Z2KNTX1t57mQl
TLvnbyS4cdyIuyMiGVKO5oTWjEti8ITLLrU7QjudNRjd8BC+AtNIF7FA0jAtvLD/wGY6JdZavF5j
ejQd4NP2nIz72LfYPfkB4gD2brbJGEslmQt5bBPtOplUDORiAEXKQHOOO5S5V6Q3nYc3VGh3uqQS
Fc1QJ6pey76KLzz6bbeuNEQXExyLuvjSN/jnWt3ZQ+9Bmy9NrPuC/rdA9n8hY0UkFR6Ucb5EfGft
2IHVQvEvwpAUIxipOxaQulVbgd2dHxu79dZhyPguJ3FQZwusWk95AhuLOOKgSucmltz9p+a7X3VP
sr09EsgK53fju8QS0OFXQeCqXl9zEUap3nNi7qGsf+xsxkKWu6ycpHC1/H9SkJD6wU7WVuG4ZpKj
GA903sqL9q1oOQGlOLgGW4FjWjT0d7r4S4Q1OWy8hMEO49K07fOeEb64n7nZPc1UlUzEmuI0sStP
WPY/dMMbEswB4bzBwY3F24JnCCSUZ0nLB/ViGqWV+UHY7OVfEcvuDDhEAUc4I9R2cxSWuaPMC3Pf
CdA8CEn3n8v0qYAmh3zULY/nSY9bdFcNABFBbDiS4W0epii68MY0/XKTn2juWbHhk+P2gAju+OKO
A0nmFyGw2YBrg06GouKEY/UaTjOLvFkux+3kd0OJeSvAAAH4/PMDHW7q1qADJ53fFbShdrg2hWcy
TXrbrBEKHlOpkTUKD8+9VwSHDaNez+Ssf2mEaOxQrhwYumKyZH0AjizCh1IDb+ckQ+7QU9gJzexs
nc9pRLxiEy3vu7FyYIkb/kSi1MSrpzI/OKAYgVzCHISQZdKJa35NlvFopvQb+XL3BDyDWe7F5zTd
CILRmRnCcweAeav8tgP2jqyCWxNhsxfytx1jtlUe9cINvP7fTX2qaKPQhOdFC2gdQ30lRQZkSqQK
HMb2ZGYJbwWfW00TjJF+1LfkEYMU8lQX5wK61GJCpZ4yx2j4C/38TqdJDqdtAHM3hpOEvdaOjRz5
F7lfdfgBJhO7iZQRgoRIglJZ1U77Lfxvla39OHnnL7PHYfH9NZjpTItGxGiika+hbVR8qut44nsJ
Oz2uFdSdsmU2w434dgMjR3bXctaMbOswY8WJAT3gxIUSPi828Femek9Kt/s3pj5ltPghvyyp58yP
zUakMdkN9eor1oRQwLsm27VCilhqcy7mh1oNjFQ6oKKKsf6JZHHoMpW1AsEraD+f5AsOIQibRUYW
+bY9Yu+jwk6uKPsPuPtVsKRP312Z1MIC01zeYy5o61egzynRhdaxr7M3CS6jXE3WRk4s+J8hxRJQ
xpyA3WvVzXF5pdVgUWCgpT6GHLTa+KzVucssfiYMKf5fS10xFQV2tn/b7JSkBWrdWBydtJ0iujI4
plHG1C3ECMMavgrLToLG7GqyJ73s29OmUJxeNFi6JII0wAGFhdFKkgSAzik6VZR3crpsQpS+KfHL
kR4/+UwhhwxkG/lRc7Iz5Kmsuzcy2zoCszCezsGwc1M8Z7tNhwpFvOJXy2GICCZSvn4jOsWq3VDC
UX/FtC2bQpWBVq8N/vyeMRqocXwgtVD6vTLeAWvh7tero2OlIOoHcfliY1hnVpooQANuOLdpIW6n
iek16CvfNBwOA7OqhgCcYvOUDCJH1Uv94dY5T4u8bGJnq/Gi9u27e0muXirXVKIRlwY1N1RIetCG
e+7mtRInt5PNPMS97teYA4mlknPFNQuq0pBOSQyLRNEN3A+Ld8c2qTid+aamJPyd5+gZqKM8C7Fw
AyHdNaokLLJIWxuJF0hrRXgfcbAQ51jy8JZbR9ZDo8AGyyk/UYZLV3TtQcTplnXzabEUGqLvIMuo
maOLzk+ugAq/D+BX/qyHFx7AOy5xi3Paf3Nontlx+XJXonu7R+Y9vtRR6U6KqfX4BF+xeBhbr+2v
4SccypESw1gxhj6CmdYjcJlnx/jmKlThu3KpMuYwIp/rirXKql5KA+ixLj9Yv6qt3736AseA3wzv
5dmpgr4tqcmnCNtIxPJR1A1PFfQ+ZhxEocvYsBOJodVKvl8WPufo0MSAzurvll9EGCvTydp2L3tL
PtQ6Nwv1DTQAx+rsAaWrm+6F/3PTCazR4odz/6FCWFYzMBpPjajbIrcrottMvr7AvXmL0BbbyH42
h/jsVHsroTQcQ4L31gN4pvq3vRRDopqVNbwUABfxScZMt0QnDtDqg/VPso0cGQsvxyeX7qMMUf87
m9xjBiW7FMPMtaQ8u6/dgURJ7VDgsJRnruCj/Yox7C3DZfQ02ucQswMA3RhTf5/Clk0ZErgCcOfB
CqMDyGyN+8OV79UqIS3MXdcqUvWdUNL1VFIlyPMylFKKu1TNppfjMx2coYr2xbK7xv3C+lhgAyJs
tm7wqwwYaso6wNXHPm7Wks2+yoK29KKCscgIvorFx9lxioqRIg99bVc72FvPC5X2mMj2+P05AeRc
i1iJkzkhazRaTScGE2HCif5QApWtGXx0QwYl/eBaoJ+9aonDEOpejVOQehJcj/K89aXNoc0mGebD
O6e6Sfpzy3FOov7aRsPr46wixEgRSBNNg8fwFUuEJTio3QrcXCuzzt7Lz6WEHZS0VwO3KjgUGWLZ
M+6Jg5W7MOXOAq5osX6PP6R1KXgtvgGt7mLjaPyaxIx7l4UWchYJPf4t2RrDBggFeE+to6OIwhJm
qoVb/yX/uxvUqHcv4lV92C+1Mya9SIeWmIKb0k0URPQ1MEo63gn/MpA7kH6PESFw7pTGC4jURY4o
OPZ3NRW3XEdr+IpZL3x7Rb/DUPaI+OrJxvzck0krfzBk5JrCPYs6ezkJQ6iETGi+4W7OtjGKj1vu
WDpDpOplsE3dv+qz7d+WRUVlYL57MRfYV7QeItQOlYMzmPOndtSYmxtvyaj8z8MS/0aHcYko6oxq
J34DpvGenf5yza+rlfl0tui6kNjZOn78n9iX/T5Axn5Mw3VVe8g0I1rDMbBkeXg1RVABDwmEHYau
w1/HR4Zs5EILcpepk4aoXS5CB6I9v/J+jT3Fo/mpzGFXSRKa78iwB0ENLLgZhzPnimqr3VWiCux5
ivdLC4CxHRpLKRmXZzcfcCA5Ljbu7FuoufjZUV/7YOJOffpb2aorkutxcxqN0dGd1FaeqpDw4qjK
DBKLg/V2XTsKccxsiwC6+F3e3EcQEyB9P6MzohnsrpPfuIkOmgXuNYIrvjCVniXlgn0yHNnk5Cx3
aVgzjNGsYlgoSZKexl8sKixWe5eS418qQaN+ZoUeGSfluV1aiDfnPAopku533GgN6KPAaL+d+xJB
wvNaPMwp6bsBV1EyH4YfWvF+CJZgEGPVfe6oJ3sTyA0TznlCjDqVcpMpc6IbfrTBWWmGgE1gxFXR
bpO+iHZVDaWKcy4ckFeZJil4TEnwhs3cG4NuqDgiHv3Norn/r6yq91HKl3ZyHxgOu+XpQZGkt26v
vzIdFeXhky/u8UhESv9mBqQw+TJbq1H7r7SRD83NALVS9l/loIquxe658Pl6ZfclkjdFRVX99bD9
JKqkar7GIO1YRonYH6P8GUUXrmipjUop/7FH55IyUErWjnpXTv+5yFoqVQH5j9HYM/gh1wQTE56d
kB09nvP7E9Jd5qHi9pnrHB6t1Nn1syIqTcgt8YtbUmqLcKnXotcYRpImIIXsKBDiboIvs5wrdRLy
XJFPu9XG/eN5DHWyjpchiktsfUyARW6xDiwwsmBB89/hjyJXr78fZuipSO0sjl+o1oMx3JWl39jL
F7PpC7kJlIcb7q8iMHKGpwk+qu+8ZHlnI0YusFhxYuxtdJ7emcMFM7j5XQ3c3+Z9fJYhbnd8Br3L
7+Id1BmHwy8wK2X4KrzIEctG6ief2Vn9Lf3FYUlpntDSc7IIJmYkcqpPCl5xEhrop0GhP/wJUWhq
m0e2btnnUnjEZsbjCvwxCb3/OflQJSkeleEOgcss7Q++0obTHtZ7nxJBHP/iHGcsGeRr8FmPxp4t
XHhwVA87GI76HCLyK9wJeDWipQGg4Ied8JnDhBOpX/FDG1E6KeiiAGviTHCcDaGcvRF0MS9gboQu
i/JYH84L49KZ7tK1mTOxeo3LIWGKuhfsumjduohFIlraqOJk4IqfFmQsKeKDMnSAuEELEB8XLmme
+zx4kB/C5qnHQjzSD571snl0/uHmctUMFz5jPE7rRp4/TdhPb2j+SPnNNlaelmOiSgc72Pg6jvL+
QwEjX25tFkj2dOURBKQHNUETuq9emqTxMGkSSzLBL99LRqVbhcW/Layg+TDsV2AB1WQFCy07uO90
oFtO6bnTj7DMLA91tdcNo36zDYgEdOyH8YQOVDpwu+WeY+P2UzbOuNEzeGOQDMyraG8SXOS8bHKn
JhMs79WcflApg0KfOpQ9PZFy8vqhg+cLzqsymoQ8M9zd0Tx55uYWT90UXunu00cxoFUWdeeJc3Kr
hwxoyPxT7wuOOThk2oWvFyYhYil89AGwUMiB8kTAtJdSivlTlALuzzfemyKuMiBUt9Zv93aXqNAQ
Z1BkewlVn57OJs3Nrov4tDZvk8ETwl3LViKKbqEcyyEkTEYE7hCYcqsXxRSpO/esU8xKmZt3dgeq
b9rjjM9Ljaq+flL6iR4k+XfoyS6EE1IOHHXvM7o7/XvPJxnUCQYSHhozswSCWweVD0mm7p4KvVEI
4mLR27t5gcf0VquPYdPRzJD1NV1bLQj04YgrVhYYxrh3I5dXA7q7ti3Td7QYmbwagmtaiDNIMVVC
odzYxL4jiFbrpp6gOenTGeUOn5rudsgogdF+E9g+BgNteot9uadmFUhV8dXFqD/Gn9J5PBeEDnaI
mFrOL1SsSfie91qhs83Pkl4Q/UZ9IOyH8Qymaou+pYEbmr0O4gqp/PQIMp8vUZNxcv0qZSlves5g
NhepZLNyHTEEI+EzjyoMeESJEUeDW52d9yYwZ4al2mkarCor94vIqCJ770lMA+6+zKGOAzUlq0FD
CDJBNr4c9YSb910IfxgRuH4R9iHNGlq2M72slY//CxjuEqm44Qeky/b86KOufP6xY2zOvRy/TxgD
tnSuvdj3gRxBzOvbekQRX+d6XjnNTSMc7Kvg4UK2tcRra8Ta0zTBH+YVxkwvET5iEa9+gCTZXpUk
B+bDK6strcoGYgi/yIUswvoA6591+C0QPhy4drZr+seJD6gmugPg5qscmTkdXveVy6u9jT6zrzr5
JLiQd4Zbb7+KnkpVWl/tl2dthVWh+D0tux8mnOurhMfbx7gVKysTRKSVREia3JBT3lhIJyY/KgBV
n5i8mu/cvWpw5LUF0gnDhddpd4y7YojeqgPtqF6H6qhHQlNX8AOvxSMtLtsYtAP8pRn+yfzO43XX
TSyOkn3/bgQZGN8RiWvJncltubS3Ry3nbB286MvN+haZth6xP0o2Va5vtXCxP+rssoI9itaWdLWV
Z/VBTSEyYma/yIfQiGGKQa+IAw8RgflcSn5CxsR/j1FI9lA05SokwYPzyF9YTl7i9Qh/ekckofLy
m0E8rKUmfkgNOFzNNni5sNmlH2gBy2iopJBUx9GCHHsF/3Fjp92NkK3P/bCWOmHw21g3zcvQwXlv
sG3BzLXYx+qGoP4wKOONf2I2fCjgAQRYomKMOyH1CtFsZfqKaBY6FActfoPb4lsU5DkKgGi6L4B5
edWi6NVRFuno0p5RTmijrdy2JUW/5O2WYsG7/jSJ5m9bHtvX7hrYVAptj2dg9rflPtGJsK/8UGP1
Sl4UxSV53h5ZBvvoHB9/FG0Boliq2eFeyZJlrpJlbfwiY53pMUR9dokaZIPPRB4Hfqtt24ae0fC2
7F7o/CtGjlFzHvvPfs2lW+OMouop0Sw/4kBA258ssdThnQZFXjt3mibyaPhlnFd7kyx/l9ucWYOO
zCIxpnypaCA11x4uA3YpZlUwmh67txX3rGuLSBrvw4XICO5UPiTWbe3cYuBzu/RVbRN1O3Y6s/rV
hvY/WsjBssVlKAxbEdpW37cZ+XrkJw2f/RlmocnKsM551RbVvzI8g03Is1V0+HFekLCNCSlJvGc+
QSlrjT3GHjYGbdUzFsN1lqEoUUpjqVVbMB1qSBcKuC5J55a9dNrjqJPe6llsE5PGLj9675Lk149U
k+1YCrwG164GeahaP09rYYzJF2FurAO4oLN+SB9qQ0fHdpSSqHeouqiCZIgYlRAc0ZKf2R0Pi2nM
eI7lW7gESGTOvfyIQvb9jLPfHMtxqDbFmUJlFCNtk8/gRwk5XmNhbHN4huJqbQJsaJXXREEs5LXN
S5fKVr9kUij8SWddk6l8Itp7OSFr8XkjdW2/wgQhrmGENv+Ou/0xdfbpVKJA/Csg5Zsb0L+esT2M
P1QdRZiz2BE7Y+A6/piXhmth3AWxwD7zae/dt67CtVCXPcmRYtW1lQPVUVMrWrta4MtxFor8MN+J
7FRjP+c4aaAlt3AkfFDPkSbG55iZ/gKbfkRWM+2mVHQFAOoGcMrHC8fBDGwMUOiMJBkkTTOWHpvI
brs2CBGKp5cRFAsE7g1uv7O9t67HuRmypNTOMdN3ubJxKqj988sweZjfnTjyWiLRJ8iPRZPlCprk
9hhTymV97YoiOoxXA18w6VrHsDU6sf8JNqRV2h9b4TYs0e0UgqqYKnBHnFZ5Uu3fWf1hdIQSsilo
Epte7K/APJ3ua/z2HjcMs5tYEc3OTCF7ImdhtnIbexBbZjlW+EkcBKf6HHY8rL47dvXT71/+KsjT
qXCEirCcflOVgGnPiM7JO9mK23IEvqNHkJtTuD/fV4rnj0xbxU0E7lgOBw3MLfRBvxzwkhiAZIz6
g1S+erAzgruxDrbaHkJfIu6U7y3kWlU8uShps0gbiNJSD8szEg3kj/pUCJPbzRCZjB36Wiu85ZlG
OZPUwGEsZ2SqhHZ5prB7TcinrRfl+DUQR8dtlPxuqHwM9EnLgp6WKAKeolNhPNzVswDLtPZLOu1X
B5qCfHG4S00PzMKsqCib+a9SMqyQZVw8ozlSUNKWs4xRzl2S5ZNTcUdxKWNjKiUB5ENrDOmMGRea
ILjl7b0nl0JL25LswhrI248nIRe1q6mWr3wQw7Ar7XQfSRH1CW1JfazDXZyY9Escp/tjqSmGkN8a
xD2CHkWpveeqLWKBzFtM1Tj4QUy2zF80C/uP777MZvSj/rgmx8W1fB11YHVvriHA7usOhyYxiAFp
BMea1ndkVrvCnsTf33vegS3yNmV29XsD2scWD9GgRF0sQC5Il9fzjG79Up4d49e7sg9ayst87Vc9
SZYfy/c4TCUPZYcpMOBUAgJ/HDhoMmfHLXnfebGykqVBMfddZKtVRzgh3PctOT6hBl5rUkGXMHoL
u87Qw6PYASVGk5tFjMrZByTJa8/Qh5AvxqUkvg433Q2dyO82xcXtbfK/ALKZ15X/y83Mb1RBFUgQ
0Jfstp1AjKz78eZs2hI/cM1coMM8KOzNYSUua7Mq9wnXak+OdHmXmB7UUvnqGkc1A7Lw2UCeEs99
lWzBzfqv0VIXQ2/8hu/8cWooSUhbBHHyxd0rONgu3PJLdr+KrmplxCDB2/K7F0B30pU1R5s0tYqj
1XHk9/141bz1rVcqIw7qSb+8UYIDkS4p33bRmKkD3HZLo5ko/w2l4mRwgu27TA8g3BuohCJyP3I1
OhTVqm9V9SUJzfSBv0ZD369gdq++HoYnTxCcG0aSiykxS2MEJP+oHd/RjAsAR6xwvQ6VQqRDnxJk
t4T1sVr8m7nRaJHV72F2KeYNURi6XVeKVsWMXLOZSs0qHqgpj3ZXUm5BnJlLFW5bbFWwFUFAwmUU
CYn1uPlSZ0oA4KwwByORpQK1dMDvS/oc0zYHGUFgtqOGI4vYOmqQ+UhrT3ofOqkjY7FsUtDGcDeg
MMcogvmCc8KBOeqAff1LLnz+8xhKzorA9+3UlWLwK/nyJuP28wpmuVFkMoLrjFlnTqhBc9DVsoCW
/PXsk6vrWKr22bQRMBCd0Ye6X7kvx9vQHZgc3QOUemwAd3ZhwqXrQ8HmeEHgNsdrrPuamz7YcfWI
zTleX9JBcgM/cu42oYL0i1D182/1Veawr4C2cEFDxJ8iEGdaaYf6+CXDSoaR3uTZsabUdUoI1O3W
Hb3QQxN0z+6j39HPG0rwVdwu+d95+CN9RHRG9Fq3kUASEAEU2yelxgTpJEteiSysFcjfL/WRRTyt
aujhVHOMd5PhCO1hOcw7z3ely9iVP48zN/MG61HzvyEurK/dQAYuxCU6e+ciQrTCixv90qFeRsv1
vyDJ/hoEsmBNtqB433B0sAd/HsCaPzxBkvxzXKE5WI5udQdadBDXLCwtK9ksjGThFQcwt2VA1Tox
wgJXoiCgW22TaaFQkAiOqYjdiGHlCglGVwPhQuwAXGMdHPLEefG+amZIh/ZZ/wYXx56ZokgPCFM/
sasH4sS4FPRxxGXI8I80NlDd1b49c9D4GvrdwHuwpflXhX4PoNwGmbK7lWu7mEFBJQKPcUyaQ8fz
4jc0KadpFhJp7wZNgVdba6HOMpEX/y3+aPzFUTANyPMnujnrY6CWvzAZWI7giE8O4wVZvb0l3cAp
dQ4HHfJ0G1z22aRrSDs1Q7VH6tIW6R1O6PscAlqRHkGOae4rDWIFxDcQFNNZX1JHJ0kBEQbcRTNC
pednF+XZJ4PFJJBpa5vY8dJmzF06F9kulETr57ekD1qQsewEOJ7hYW71oOuSuObfaWCUHXgZ5D3o
QHGjmmnNDFGe9VeKPFa35bdATWplSYxv8aG6gtRoTyGYRnFoUcSyz2U1sIYxHUv3XPFrOlO6qfHb
jd/MYIZ/KhNvwDSod1HVwlkT1uWBFDBqiTNm/xji9Lj5CioI64bNnp3P9lagybN4xzh5PXJU9GDu
XGqHDzT/EO/f4KqJASVfD/p1Zdg492bSiPNrtAhH9X4CkHqllcHC08HIUR5E516fF2fMJGJLF4Hc
olLTVZDiVYCzmbAygifsp7+WH6IjiiMroQD4woaDiuz6OmPP6cw9aSl73LJLsPcNtHFV0yb2/2le
oRzoh53ZcmaZ3vhT0hDklm6o0MFwqSZPqs6F0FzjcC3ziKUpZ7GoSbO/aS2G9mTTx2hrbd9uZgWX
H5cxas21WBMh0lSgzJ/qifOvkRSx2jGTorzzfcQfZYJ9NEWW5scwlYxtnZ4+wOo2wiaa91sgaEz2
ivRY6fBr8jXCKNaQRRMTsU0CHti7gnLzXHywvFai6Ndmm2lw0CuuDWdhK+iZH/u33qxAaZsMcm40
0Xf5sQrSf4+4eAQFjTRkXHlAKBQO1G1lHjtaJVjWzj9LIVqOVCvYqmBdkI92q1xnMKPxU0Amg9lx
OfQLrDlpxOZRfxR9bVDbqP8lATmVIotIoRoXHGxAMqY5VnTtiaeTGn2sJ8focKBHKXLLH/6XU+ii
7w30FaDgTiDpr3fLUTjJxHXBFqvwGjbUYQ5SA0+4QGkHdoweA6H78X4g7HI1qhmuGb5ELd2noDbB
5m1Bk1GAPDBy9MgzhwvQALETE4fVlFpiQAngKHIAgV8OatYDuW0FC2AMINdQLJziHJr17F6hw3Xb
5GMefDa2Jq4dW0fR5ns/f5jI5VCn98TqEzFa6wifUuqRCNoBVIxfvEri46dIDii4QBf/QstLANWL
CPuu/qrEcOjgJ0G69iihLXrWG8GG554nXDirIpGCkChi6iuWnCFSP5fXzzJFOBY0jNNDok6y8EVG
l8zm14qZ+M53bO0FUlEjQEySN9KsYHhZuvCM55CKL2J5yFojw1FUzZFlzMMBng7h4h/MOVpyY37S
uBrtFBd9mqSLolQ0z5O9HFqD2GmJzW4MV8mQ1WGRnz+29h0hNRY8JItX0FZQPj+/bk8jmEI1cjQH
rqX5dw9tk5tSNrVg+x9rTnpEGEf4M/d1JhLTEGf1PrEVAVyfILqSUUqwq/AwBhmWy2FUQ+fHUyKz
I+qY9bNmkwTLBSyhl4k9AsaqeKTLJd0Pn1mWaTBSgnmJLN+8JfkaZdJ3k8Jpkf2daMckUQZtKylA
jAawvIIWd/Wdk8c3Bk+4/+HphY1tnQUcDfUocrjyYkRd9tuXlYzzK+AV7WlUvucQ30NgzHrOzehc
Kb/1ffqD83yXnFY1u4EcRlMb+cl8KZUoj7etCmMQPk/+BFrB1GxDsi1kmewXCsaeFtiTdxAo6vhV
XBorjy1sVd99U/7pMlt9f3jiU+dVtkhxSnekQFn7HzPr9FA1pqkTnI1OskRNsleYogzJYH3/h3f+
MW7fP3tu4de5Kxf9jnfz8OqIS2yw7yyN9umgYundYid+n203u805Bq28mQWDYC/Gy3Tb3AmSQr2w
ARujbBzlb6ttPx+WxYOkKro+/Mx3BtNOko7H9boIgOfRgMh969Av+WZLkPHi/862jnzAv7SklVgM
2RNGhy3eEA7tj1OZpzWWmUVe2LrNaiwDF9LArN1WdPpSBq0QPHOs1TXPPpox5NujwW2ELKBj1Pqh
q13MZbwJPmH/pWM+nNofRHcA+vVAMPRtkAM6+fvfIKTql2j2i5AFSexFndm07BH5ah3BgmFWEirR
a5u+16t79mUEzNj53YHri/JyD2jjRpMtA7u7P1TQHkAhrDvCKcpf1E2qPKbgW0dB8spWZqB771Vm
eIgryOurxCO8l4rPXDdEv51ztTghqsJVZ2OKo/uCTbArmSxB0OcLibBAcCYalOIQt1O3tae4FTxq
ApdW76pLN5gSQW9kJUtaz9BdvCkzoxWeay4YP5afLC+SveCPST+AqqjtSE5g+bm/7AXuN+zxJ4j1
ZdumT3JrQY2Vz9fstN6CatmL7G2GGGz4cuYSLz5HijEfAr+sjY0ZoALduQPKGyOhyw/6cqrgZxBJ
hP7IlTmW/97sBXC3JvkXhdfy7tD4BmIPQmg/DER/YeN5ESpwchec6XU5XWbHiYffCYtidbLXiL+M
O0kxoqmLg3ulaFN4q3c9IK1eCDUaIG+21ExrewMz4Ufl05sQB9TWZ7FpttrA9SMp4uP41DNR8t8d
qIHdIv8fSq9Iv6H+/V7T0kPmf7pVWZYLZMAKns9Z+YaijZMycIXsaoGFBMc2La2DNNTeIdY/co89
mSdAq+MSW4WwN+v7r8SGaayJEYoTdPnHymFnKYvyWDfrVPBU/cfCHyXfftl7gbXoF3uSmKkUBIMj
Fp9U1Ipwy11Ogn4t7DztDS3cYe92w/GTdJlSBjplQLSNo6q+2YB6s/gvM+a/6JX6lQpnKZriOOfg
ERquOlP+eIyT5ArBSoqSrpMjxhFOb+SprDmDfSxXSnBXlfH1qOQ40EtN4TRQeSN44v9BjiLu7Tc6
vd9qjZ22Tk2V6D8rPi7uxCHcXVstZK0FzF3EWYZuCSX0EGtwzpGldX0UHBQMzrzqmXZmXWFtpNIf
tkrPF8MEsV63capseMoN3VqOcXmgErvfSSBHXo9x94UwjatGNJTEpD1WyqF+X04TVhl5j6z+RPKd
dkaKIvChbJ51KB2OTAClfz0XkYsJkvlcv8Q/+0uH0fh9okhf+svflTwcP1SU3dusGofbiPBXOGb3
ba/2Eu45nUyK4crDfM7RAa5Qx61HCUgJb3zwd6tvZm+qTWWcMgM2n6HBgqWTxuKL+UwWT+ZJDUPo
lVSYkhIv217Qk2w7DXzl5dq07fJM0enBloimV1aymKqtsP+gv+a1LGVXqJZhRPL11ayTPUliS3dW
7T0rFA4W4Xz+dz26Fzy/bJeJymlloYPLJDXOqpW6QGc7Yf/0vFWBmacA3MCPoqg8LqjrFpiVoVJw
IkZqLi+FFGijTY4YbafqtpUVp889WeJrBdJCdQELoHmvpMHJyQJKrzB6NtPR0s4B77mfZ3FVTgCP
Gmc5KDLJf8xFvZ9P5UIiLocbYi6+kh51R1Vs8fGZbKfD9gVQSLdXaBSHtqM7DMEdd78lJmQaLVX6
pldjnqrFWl+Il5FNphNJwcMnIcJyKicjyHKk6UNHya6QxbhuGM6Zu6BMVaPu0cd19lmtdbUljOQh
cmwzvOCT+RtsNyo07oQVVPv+Ll+d70lH4QeV2T6Y1amVRmqxRhlI8GRcuHFrFM/WfisETYmWrFhw
Pdf90XeDs3LgvfMVyrt8+c2CHVx2FVxuy4xtUxoblf0m7WDjbCZNQwThjOXC2eS47xIjCsWvJFMj
SXgwcQSpxBE46oWZMdH0fkSH5M87Y+JWC6jloSBilO0+8+dk7XMDJ0/CKrRS48jgWMWZFFNhgDGF
4MZjUdA4B5IQCpbk9+dWbk3gqm3eyY1quAqHLCoIYQAADF3K8b/Q+W9rUKVvA5ZA3XWwWW4gPf3G
VnRho2VW6hJNdDE8qoOQLzX9BF9uqbuT/wJaLBBUVmCZEEioCeN8mljS8QgIjiNINcXmGRwiguJU
DGQRKh44D1ucmio+AD7ZIfEJj4YgiNiRomrlHXZ2ko/dcg9x2ZAsMyXriYYwHlthyBuH5gUs14Tk
YK8vtEGbFmUm6djtRX8e/85w3XJH1psxu8W4SbgXhvnHM6fvM2aS63HWAMf8HTSIOipifBNirK9W
kcRlc2N1HFmAr9bPwldc4U64bkTQHaf71cGKHWAvUtzwmT9sK3vwrnG8xwf0x1Crh7VIfPS5yFjb
/lUr1xPNf/zl+oppnAzuVp1M3kuli2pE+1esLoE0tjp0Xrr8TJGBvEp0IUIG8aU5fDQYEt3l8YbZ
IL9tBxz45UUOD13IT1h89jJ/clY/GbGOV2BzeeO+whxb5AFk/EnfudzTHZIbf6ulxfRVWZKAIWT1
+79MfTI0AIGXSeOI7rWF6322tcm9X+meyaVyZ/rS75LF0mnJZIiLGG8TNHAS40g+bIkzY60U+hlk
505/h0awqkqolxhNfaYoAX1dy514Xs7n2pPpmkatQM4eoZDtstCZatoHAuWUfCnEGmffNZIJ4FNT
vkUlH5R+/feUlST9JeTp3+albLhCUHDSqgK7efoZDPaOPdpsw8d90NMm0yIQr/a4Tqb+CEH8Ck91
jyHjMZbUEsjTAfIRXKNT9SwQdXyZUJBNiJ9snkmdTNA3F50l+fKNKDFD+tXby9dgdEnXZ4hoVHf3
Lso1wlIu92k/fYtxU5zPdm+l1n1WyS210dEXWUrdAJMCC9x6Mfx4fxiL84O/ZJqheC/7uLQO8J9W
0tzzkbXt8wTesx7GnDdkBG8zREv3iKLCRKQcXhi1OhgF1ZJE/KsevJbBZQmW6W9NXOgSO/mhu2Lj
REo4bgKcQGvnBhJovvupb4niKQXAKyfyoKVoU8gVySX+mqX4CnBp43wilaNXdkAL+BWuPFVrCs6K
ucegfoDvW/+pv3p9ItNwteLWQ+VjvcBnzJZDCrYVW4/PR3vgMz2f67QsJomNOPbptQuRTkXFkagd
TpZjvFHec/vUNxCvVXcuuK7xrkankrPWDVNSO4EXwLlkdP4ceP8XibElzolpg+ZBGgWAJ3nhrWN6
ACnTOUBaMZJb4LElcHPKJsvuidnU3qXYkPioMz174BIT/+n/UEhgyYploX9/meHv1Q15iQKfXJok
nYRufIfpNRAR1/NIqXzvzMp6ZSFN15QMtZomAaajjVRI5+FHpA77+E4fcXe1J13FkkmIwLn2aYd5
icmPhKsMwekZ2q3sRYtZTsUPIeVzSbSQL2jo8zePB0MM9350AE6AYxx7uGfdY9B297D1hYZrsjyu
hFTAoB51h3zHviUa7vU1hMIcW7V8WTd5jUlzo1/l3dBkIfkqJDHapFNpTXUj/SxFqgxYscCzvoyd
q1RNMojCs8+hhhrU9xKslc0UuRSlamsYeCuOFQERBxMwl8MC8Fa6R9Ru+wkXD4lXPmiSa4ItYm5i
1bj1vv+mfgXjr8o1PIOFG2yd9o8T5pLR2c5BUFTuODdrJ/XYmn1nYpRJBU8T7TmSpmYumyvTIkJC
OZjU88CctifUoehzNOm8xFdVretgbka5J4ksoZbBZrdxxN1qDyY6PPxKNoqwun0xOIoSXR9hI84J
evYnc/aLHA8nJbUJeMyTXNQGLOehxAYh63Rl3MbQW+7gQ+fHJxwwhHxAXbZTAyPbyPN19Q2XqZVa
CiZmPIcXpORXTs+WyQoQ8BsUBl5285YWI+kXGSjrtb/BZGDlsXK5DK4dHS+9D5fWNhymVFMdCiHr
Q4renB+XjGQon0kVVHirsumAxg+kLs/JMRUCAlyfaEkiMnGXrIcxYuA4ZuNVZKpvf2KMa8HVLadY
tXYri3OmBOvFanrMqWEkbu9nUGAI+qoeibhnQWwTZtuPqgjRQzYxRFqwys5zZ2WQuzwjBVyU8HOd
W22sTMII6DRdM8GtTf36L0rux/v0ouBaURT+uVCha/JSYdWuXjXjADBgv5PeccCZZ7lzEDolIFDR
RSXZVpokeHDkfPIBZ+kmFUpa8rcPqiuHDielDPqw9gdRM+avsx+YVkn0aTXCP7DwbPet/15Wj0yF
Tx7AnwqEg2UOUpsXykMCRZusG8/ekV94gEsqQexFmKDlpbRt5i3jnjap27QSl4xIYBr55aiK/248
eEZe5OUeLzOAbbEyahZKCfcjutxkIZn6Hs7C0Ut+P8NKiGzwZCnPj52cZI8oEMbDtsE/Z2yuigR3
twLezESSH7xinbSI3wLc2Tw8S6U7Nl1XkQM8x/O2f8FbK4iEPweTxVEe1ANqiiemA5Dm/RKhGT8s
u3iF7NE3XfReGj4LMeNMhUlV3H3/dEwr48ew2Miey392DgAYSyUb1pC/W2/RSEDHhpxHEYzInrxc
V1OwjbeVzZys5QfOECqxdFueRgQJbZngGBxYMTvPIev4UumHMzblAf2drZA3ozA4Q9YhRJqja07a
S0SC8ILomHYEaNiS5am7QL2bRmpVc3t2R0eaUowITYuO6MCv+yppRA9t7AKdEx8c449Fg5tQQpLO
mtj3BNONfiKBH5kJhi5nIKl/QO3v7m9fUFmQjSSfipelKGv6ZkPKrjfyVoAwh2qa8SBxGr0Lsg38
ZtE1vGzd3QOyR0/4yAMkBqlGNx3bbmkSQZND/bMGcX6nlvLNqtqTjiRTulEwWTiCFtzimIfWw/Rs
fpKXDRXQtx6hJW0/678m6urMo5k9mmqfhSBsbEJrVpa7DeQFPbeWcWJAxQdqJbVUoBpv4+MBhoge
I0OpiO0CEoK8z6ckXjTNVFWtiYvROp2z+yFATwBcvR0hSdmc6WixBcfetGRQiaZuVgJ1YwRuopho
k1ked8BAqsWZNDcJxaf+0LZS3prdAv+5pOQdp3jdFBgeaT50xM7W57RManPi0MPOzvvD0Krf5uel
UBEVOuUEUURKcRQ0oSLxAiK+CxOhbGli/iEW/Hu9i/hUvYngf7Embm9UsaQlw+SpI2osc/ZyKsgW
7QeUA8StvqvlvE5ahfp1bvpSw842mvQTwlty5onDdDcwip9/a8pXIh6NMnov/mX6YfVnIiiAE6nl
a60MOHnoOTcbuco+pA7Lx+byxyrYhkELpkDaAKf+7vUx+k91DzDzY2KMg861PsLlsBihXNV31bLD
R0EpLel94dTJta3pW7p3pr76F1IA++OeGHzLrC3XRbLtd9TzK5g6FKr6Z9YUVhPZl6SVrNZQDZWn
k5OsX/tYNJoSRr+0LMMN8zj4mQFut0fZ0BJdNRZddub7Z1agBDIFdpfeQ9LoVGBKLX2ZsVm7wUBf
h3aynDX059yZXb4ccUlYYkuqjnfG93h352Tl6WXb8Ut6DHcCL4L2r5iwuOW8x4wR+sdPui6l8oA0
WS7H2xLH4fEN3zcsdIHoFqDoCwIef5Rng9cB6X42h01TeaWU7LybtoSysBbJY+gdgv5K7cX3pZMt
1hRf7MNLjK6zyQRSSiV8g/xvGKNLgZiyimE3Mkn0LMhWcdlb/7cCFRdoyy1vW/El7Hd5YcNAnuUy
FlIqwFqWLRLQ3uNLYXV7NmQbJdhWAikW2fSnlkbH7KGgvIXzAz+2aK08HRPi6qC98aXqAmMWQab8
+7t9PdrVTIZUCpXsDt4A9KELDpuIvhlqzYYPkLApIgRx4e8VKg5/HM1qxU24IT6bdzjF1JdqCwf5
qT30XLUqnb9yNUApFHFLnmU1RR2U6/H7Dco1l4yH0ywPiYGev4dx7ZhQbfhOx8ff2xL/yXndYjoN
TQPXFQdui+ShwW3SyEMiVzZlPBNUU6vfdWlC9jlvESr61PDvPg11payVN4FfRpglElzk50H6hmCi
bN1BX+LFK5eHurIv1zA4ui85Iei5XXLTVUB7h9Aq+LybrMGypzm36AjSZttbPlxkxetrXvSwGwvR
eyCt502P9A+LYBSQYUprHOyKMyk2s2f7T96PZa3za7Ti28+cLY3o2piY0zq7vHAamuiSJwR/PP2Q
nBd1BYSxJelJ3ZZmzmNZHSLxGnXdWtWttpehpyyDOgQyvvgnFFLLpqXUPOtAjiW+Fzw/N5mnOu3q
5sdrzHiCEGMxuVBPk46OUUht2mBnqML6pI7+ivePejLpGeJqROa5UtCfoAo9fBDhjLw5cEZNqi8f
vo0kJ0ueVt+0UOlr9co9tEac+qt7ClrZLwV/y+RpwsF66FZ6aFNorqNpf2lh8sALbzJ+YTehnDO1
5gMIdxNn5fORMbNMC15j9l0pXgiUtVG1bkYWp7S/Pvc5T4H0vGEEfXlqXhb+1K4N5ZgGryaZO88b
irfEYrCktTyS/a25LPxECBdaV9kUrByIzOhj2qKq0eB90iOod+hr0JjA61pkvpBVR0/YMd5DfWax
vyX3Dm4jhZDKMPAD3pujDQnhAJwLIYIslRCBZIFGTJDrut8KCKhNdBgDmabIeXyhxVMR4RRpJmIg
0gNZl/lHucn+EjCaEek6qKcB8EHW3TwDlZD/mt1BSNjsQzrMYmBke8GDklhEz4Ooh8ke/dJsPdsV
FTnnvp/GdPjX0Uy8Dte3wCG9eVWY/o4GL3J82T75x/JZG1nXMNNzIi5J+HD6PIhXpjO0SFgeqPIn
y83pQJr+pAH0F5tfcI8vC37Dyh1nQj+DXbp5OErW3f0EuYuxKf/uzMr7pPQQHceqSddfUXTsYjf7
y9bXq/+tLTn/CtoZNO3kaluLcuK0b4SSklYwDute+RM02rUs/HkYX5ejXLBCTTBI/NQdTMoBytOA
aJ+h1rMBjYzh3Pat+Ik7QOMGVjxqcRlXDdKAuCLMiH/RnPuigu6AkT9KOC4C0lbIliAeLq2kB8jg
vS8XrWilKRx+HJS1yNU3kp4Ss70Dl4OrCokb1LX2Mf+i3nGw7/lEVisO+5r7fYDMnq05mk59GRcH
6zFW429Z+A3exqvpIrZt41CmUAFosg2FVVruipeIsxjieeugcSvMtyouklO96mnnYVZkmQ09VxfK
A0brglEA6R2gAgiZQ16WmA+TqXLGUMX2UtPOhg3KaWtGrMFH1KAJzCt9JMwtBV8payklq/6ojSxD
hJLmRASRxcpApzLnZf48OumSdX3YNKzGLbj7fFuXK2VmTlHfnSbZkVBE+mXZVvs29+wGwWt68yuY
f7qL+GntBy+hXVa8nuAZ6fF0R4ahH4kcX5jXgZ6OnZnoVIiswcPDLiAuAk9CbN1KIZ8/s9BMEMgk
mMNjo/5ujL4fmbbpVWr9C3NGqdxQv30Vb9E/pn4J/qFlwGizwNpFJG0+L7jCMsAPoZMwA9BJhD9G
oY0Wkn/gHitIevorXMimUuUMalOrQGfjAjdMlAgkPbmVTt5ARHX1CDwpipAKOm6ZujQ+fy2XZHyT
hTAzKACjKKvgWAYcJtcCuINhgiJcCehd+MwwJfsnLcAyGlncnGueO3w7KvxPgtDCHLf7tQXrI401
CtXgDRkliFVhzrGhHVNGgRYo33bIVMoF2HNmbQ3sG971rcJxJl6y9dQydJAm1pZ4/8dQmMa2OAsN
+K0ulCv7w8u2k/KXM4LEZG4vvagR1zYI1T6fIbTbh1PdMMmhhfkCCUMU16BWGpcUeYxFSfuGhpIK
6eR92qcXQw4EzGY4BYubJ3VGjAezQIvf6mztVSBmMYog27o3o+IqQ+fmS9yb29y3JKkQtK3QwCOd
2I+4/Ujvr285JOKD4REu1r97SnfH3x2zSH7WYx7LXQEDKMCmKdHwgm10uHnZhV1rxKpCIUWt2rzU
M80YuHlLGeW9tOPxSsREnewrTHBiNaoudF5utYo7cv+wxa5yE0HS27Ios7iGWjVm4wGQO95Ohp//
d2lu57/2/tjYYSgyOjTwDeW6ESJRytJYtF++W0+y5MVCqVh016RT8L5/tGZnZ7WzYqMhtr6um58N
Cb87uTLDpu7i41ALDkSfDc/8zGzKzdXLnXDTY676nWEuFC4WfEWvd0BERuvAiz7fsxEQI/Je47+B
4vPA9zua+7u0P97g/z+iwI4nW7DD3Jg5X8YcqvxXgOOd9qEpAPFbEz89246O3j5knb2jr2RHimI9
uvr33cIKXB8Mu0/T+uvKGLU98xplWnxQnCnWVP2n9kbMj7N2AoH5Kjjb0b1iV7Eg//76z4EGv0j/
rf6TeBWXURaU8PuZldPg1ZCY2tceLI5q2KpW8lDQQYvOoi2AvwGmV8rBe595UsMFvgGlXy63m9b0
+vBVeLl6AgmjAfK16WuNg2ZCEFaizgbUiKTecUkO2s7CDIE506A+OP8Ab3LTF2TniQqm5dx+Xppx
rwLth1rCUDckZlF1rlfJQEqf8XbesUaNMEvgi6eZpnPul7GsdKcJkcDHdxSqQ/pfX0pTQw4SBxDa
9TBTNRFHf22hQ8rzD7uouNk9AwNxciBVjHP+g/Dse7exfK216SFJelkQwR9i72ZB4UfYcJEtnN+T
rB7pr9jDaUuztw+LXC/qYAhlfaQ9r2ydZiqIbpHw/xJ2DTjdsyb61EQXumXeo5xqvYxGbpe5r9ug
C7cNcdsN9SkkIQofV75XaSD8LsqwkfW7G9YSHw6KEqtfDvZijObiUtGVr34s93M9m6BwIxEqGXOf
Y+elds4S97d5qlyIMAZvN+yyvx0MwFKZoibk9rQsmqm/QhuINhMgIevxmwXHMc4W06xkZWXnYXvi
IqV34yPfdM+qPa8ddtXu1oZR5B36LYny3mFBv6g1J/ffedaMcRofZF0ARRIcDPRGZhokBm/SuccP
umMALrUg74W6+Ov3b5wyJIli0NkQ87BHlxpQv18Q1In64RuTlSAAXaJsBTKZhKNAEUssfPYqyJU/
rCoWy2NUIsXQvNjXLct2drYHOrS56IkE/h/SlC/tDA28bdr8nfzqa+Weq+wx/nGyz0lsre/+3zWU
Udt2PCsx9Bvu+2LMUul7tl8o/aogbaq4SXxPfpY5Tmq3kWqYJKhEVJqQoF9mKVfcXVvXqZaB9VqJ
bmUMSHad1nwpwZKGmX5xo8BigHWjLcfAtosnsAxwrcRkF9/YU8KH9IZYlS5mh9XJjv02YnUaSnRm
qKZzPgRYBpc8fY+Jo/9F6YI+5A30fBqUsHlqqfiPsJJ2TeOQh9z4tZqfRNBltEtIXKQjCofd+ScI
Nv2vRLc2vYvjBPDMyojS7gKSF7XTE4MUKD1WtDUgnLjvVI9T8YW5kcbYgL/Tl1aotl+HmWgldFuN
67hMUta46Hjj1VQeNsNI18UetmF6TAq6iTf9hTyURcsuUmC3msp7WfB5x4YrRAkuzHT0sxA5b2X7
Pb3sEk/3S1XiXPuTzeF1Z7KaEZaXTonnjIP8KY8qxRTm30uyhJS3o6vrLevhTuasmyT43VyxK3lp
H0W0SQS5v90QlCPt6j6eKRe2I1q/QCmazrmHk8weq/z40US63tVQKUZ3IxCAPxmZ7g/a1Ml7GClc
x931lkmwiOmkV5S0XWROVWNhxtObgFzA8qHuYza+P85HOXbwV9HtJYPRlX7TbShaafIy0LDeK2KX
Ua+4U+r11HdH798I+B5ZqUAEPv+m6gd1CFwurcm1ieUIH5tmP32IVFTBUkhZUes88AjLz9EhgiCW
3iRHUpJp8kKyl+ayiSTD8hMBMqtN0PmJ5qL3zDarMj+26VJpFTSN7NER8GkcgtoKlLqAWWT9vpcB
BOc5At5QhSNWGi5VeMY2rU57x8jQ0ZVRjYwRO8sbnw+0ipp+yos5eAKsnEdA24bTkhDe6MiZEU92
we8DoBi8aXs2bl6UxpEvO3yM636oNeNjhP0RyNc9LyW0DHRdjrf866rTUS+5yoFnaM5/W5UizYjJ
fgQzSiVgYSDBjirh3F8p5iIbb1AzuaGaUmaepBaiGzTDOCfb30YomhAn/Hdmfgqg3broJIS8EBQI
K3ewAW7ejKQTIWT2OPBJyemYn+uAA6PPIs97Am7zx/TXJLoLoAB/nQWW4Qe4rjEDbHDS9VgfYtVh
YR4GF2UoOBwGKAP5kGzfMgrPTgZQCN2UQpjrt3/KZzEh8OGVQnq/KnyMdOQgptMnm74VKyA/Ykbs
brS06LTQgKKl67LtRW3U8Sv3mVOWc4EWuEE/EdzFIBU6r/AJAL0PQkkJ+MfXivkUt5egg1+A5ohZ
pe+l7Evh7Vmz0s/MlBZBwFwvjEhMHEqWaidHTASHDvyYWukTHUZxDsNlNPpw8tEU4J7SsrT8ncsG
KIu1pKVGVTlnYS8g18E/l8ODB6PjTthW5znK5ACg+oTsV0NcdmFbIhC3uf6LFQ9Jcv7+N4OkgK5r
sqfnsrAAZRQjIFgyAIFo60TcIxRv25Ho4YgwFqKQJhRCQeWAmt+Boco/hs8fJCPIcbFMQTuzqV8Z
uL3IHO3/5LWf/4dkKy6Hwl+HOuiK3+Tr6NWbRKStQIKNYZ6hdTTua+6/CILGkaWsAwrjQZIWNGRI
fyc6vxV0+8+pHzasazb2sw3B6y70LE+yrDZHeLc+X4kou4gucJe/R+j+ui1YEOx7JbNJH4Ox0UT4
lfKBck2Az5Saae1UUwKLNeat7/I5qdjv6WgWqKCfUYWt6G4P/zcLaZ/a/fZgkSmT17Gwg+0Pnqz+
R3k6WPtGg2JJAsI5tlObZcl79+wGdfDr8gy82AXKUoCtRcDRVi+3U29EP+T5XPkXTQ2ZMJGkWrii
5+Jm1hBQvacEMgjvX/Ojqfg1KV73YAbpwSqgYacZ12oh6/uWDjWeV8XI7FAPezSnE6pK3P4t21Z8
m0JH3Px2dC8sZXCOx8+ISjq4ilZklbTC1jRoYQZlwcaiTBY+ZRGng2rH6nxSz/efOB2w9H1HTGjL
9Nk6SDACRQw4V/wbgukjvw6HwrhKdz6O4rNkjd+4jLOqveMUOXEpElox99ZhcobXCM/0HP5/3LNT
ImEln5sJohADRWgOYiaI++lEQIT5RZQiyPkikx2Y5QUn4CZbjjfgtKe35K+VF3xPnrxpR7ItSlhm
iPIVUh/HcxIRSmnf2ibifucLIGWYjvt7nax3OoIRQ/pX/B+eAIJAOrZu8C33Zk+O3gMlDL57iJ2W
xw33AUcUyFv5ILRYfR2hwfnJjEUz6uu5sd2WW+03Vt9HnlzX5YLFU4Lx6Rg+9XT2Xmc9A0aziqf8
xLYBsOplkL1pQ0mkHtuoJyOWQz1KXmLIAKtQaWi9jGP76a4QczE6QIwN/d+MUaDXfiT8vrmRmmJO
wtIzued/vzuNgtWCxmMrR2O4g6U+a6VnU2KppRRyg/MkBy3NNiVn9Zf/p7/q0aDOxN2RISWFSwsm
t0sUzVttWtEit5ZKGeae3euzc+ToYVg6nvgOGBQd6ymXFuzpcsBgvCJDh/Teffc37GwAtb/7Ro/i
dP87lN7lp+q1N2Rtav9rCJW3Qh8VrZr73/MzDlYX1qH/AM9v+9p9nQuS+z9BldJwQA6lquSzZdxc
IPWjF11GdCO7ntPZqG7/xqsNwH4GdVipFAxioG5hBT/PT1tZjiZOJ+5GmVtSN9qn010elqMOq/sP
EjRIGsSuJA3PRUvnfKwwUADzv1IyV67TyM+ULdqoFb5K5XIcilngYkp/bfJbj5wHDIgXxcEeSiUC
Yy9Z0K7mAa8zRTZswCVYEjiZ61Y39VviWbpvfrMRvSe3wLbu3wkaR8mfhlvPOD8nHhq3DpKGvV4c
5J1fwyVb8wiN2yEWhcjF3vbcQ5eZ1+9i1CzR+jnKYGeuwCpcUSmskK9Ipz3kXXq8FJBLKaBPv08d
j/Q3kFtptTbrPyHx8iEeFqKJrA7A4vC2dgZukT8nu5UclRKNukX1DHgYHEh/t4qUhow29SAr/gmF
MOKevMfHdkaYn5Dqf/7rY6mvkSStS+WZGirvAR+aPeL+c2Udd9509JKMgUYvsE/XPR4mw3Annfv8
ocAYfQGKk0XHAv80YUPytj8lt9BHg2NUROZVkI9CLoZkydjXJmIBUONMwOca74Aru3HiYqtR6wkU
uASSyLmir92DWZEKrac33zUPYeP5mxDAV0ER7HmGZc+QZjFitTtZ/rw4VTzvuPQjE/n69vgNXGyh
sgMW9Vwf57XJzJl3YniU1oBaO2oLwfJlrNvYUVwM5syX7tt4My79XX5rJ/UVP74weNZx6DGyF94d
iFrMqOsWj5ZoIdJ6k56nypg8WINH2ll5Dw+pWFZ4yI1VGCKuNQhBlVnSKrmg3vFKjjHAQ7Lc4htS
3QZ1PiH8pQFaGGU31DkQ1KAHl9kdQ6Fo5o35lrTDUx5mlgcbWmP1GxbKPPN3VxLAJNs1nGoGY+lv
x9x0QfrumB9Y8Io7kSPpQ+buHWks0+MTPlcWd9YoSklAHbhyMMSve7FyYfkrTTD3NH44fkpyQo3a
TSij+NMxXOvIjn7dkGizWTAS/Bb8EGMAoFH2YC7OjWK/07e6Dv3NisTyLzTJbiOuvPC2XlD2AOQ6
E5C/OfVxxb1YyRNa6rqsSGNdIyTtGVJpojDMQu+zSdFNj/j/Cv4RN7gQdJUAYtmkt+7ZjrqjXquP
JdiYoJ7MAlU085IPSPNgrhyz40J1iqZ5o4acrDmPL2MZWWuj9vAhtEbMLTUqVCKDY1aYuvRJkROj
acR3esz3/Cix7Af6vKtSfaYFVxxR/Ig8qDPS55QFmpBadTf9mncMvxeqzsAW1hk45NsCgP263MmU
f48hWkjJJz3D9AvCgmExpSo03Ow8pwkIl7qioy4u9R4vi9pFy07eghp22xaCvpMipNh+7bdY3r4Q
oX49aaXlkFGdeNdR1K22HOLO9kxXz/78w7ym5uB2KHj7Kg79XQowy7uNadNV7EnUSDxc1K4DJ6ZQ
UF3St6fxrw+75tOPYDlk/0SP6iG/yWCAwjcdTcWO4+Nkrboq12ESO55ROKuzQ0LRoCdE8zj2QDSm
NP1MOnePb7v6VbybFoGTZkKw+7lBKYubx45cJrHivin52Pr+4ukg8nGBnyqKaT/vq4bx4Jk27rL5
j1YC+jW9jkwQBeMB2ucWjTRmiF8IHa1pH4OEd6N/A8U4dDPvxXM5Ca5MADL4fhC3dyTe9zS31ame
XlZEWF2pOkAumi3HlkXunDHAAIcdcT2qSyFCDPoX6HeD3i5IeEUSKHadGfk+9t4eZhCKGcO5++J6
EjBTZbS13G0Oi83Tst8McBjyyjnXfbMwM5vfJeHseGGSHN8J1KdkhNoHVO/a2XJ9xtr4AwufCQXo
Hj2WfJhIicpB2ws5+lenWwAO+18JlnNoSziJ3nXWHpEunql+eEMSHGUOrAEm1UqM9oxyqtbHe3sV
a8tWJMT6z1aJYCjB+UYZzNvIh6Vhouz5E4ZBi4Zhw/dn4JbABjYw8a6PWv/FfM0MwdoMvEUV3Xd2
hvRl9lJTz5G1Hg0j9GrSfyoXCTydjO/efHPRuWVpSx339fszqaAGHsuspj123GroGpc3DI4VMLR4
E0WRqMmvBqKhbcTYVGZ18quHtEJyTqF3zlMf1/U98x0gnuon3kWg2wkYBCDTJ5I9uFl1FbCCxcmV
lWyK9uA4ty0pPmc41HSFPp5jzMOu9BMIoAWPTRYhcHTD1nbEIZNc3bDPUwJSHFTkqiCw3CGbDNuv
X1EPCaobnig9PbrWdxv2KoGKWMY5ui/MNk36UIWKYKzCG4tGWpjlZyxzbI3R1Wn2cWMpCNbZGOZ8
XugOTQjwwPLKop2ZEne6joiKw+t4+DfVqe31Y8ofMSbMy1sUZARsEysG2rFRFJO2aa1zED+u2YSS
Ozzd3QTPySUR9bxoV1F5W0E6HMsecwRhO44D1YsB4cF0LJfwoe9SfO8vZY7bVLs72s0BDcGTUIOC
9yhxlUeUepPRzIJo7kiJhInYOuM+Zmz+ri9dDVLAB8ZNdYsnfRVKIGyNnP1cBrscR+jMFqzOXwX6
EWk5/bEozo/o/0HI0XgF/LLV1eLVW50y7DGlOF10U+qxj1kTWJQceyT1vhhuhJ1hKcVwoxGAJguN
6cpZ09mm7DDabOKVvqvG4E1Zs8GzUKEYQbk2+C7ucgfMQwa1v+ArOX9vSQfPxHYTIRVnYy2VIBdb
0ZnrhA1Pnx9F3PcoEtEKgIuCqdW1rIJBOzYP8xqvdIpFeTE7Ay/REFsrTUwENWiLu8z8RGW0Racb
7zQL/LtFjcg7PFJJSf4SPCP6d3jBJ41URBYzuWQqhuuWFDxWiJdxAb0R8+qfJjGalBvO1HWT2Ugn
SavgRvcaqhopxukw8gI5wRtrgyhFsI7/uyu10cL0DtD/HMI4DxdMoE3qm+PtTLthQFSaupS7WO+O
+O4GptJ7UuMNpQjBDJDDzljEZ/16T42Fz3j9H+veThR49m04ABio47sX9GKTvFFuFX6BY3zP+p8r
UVwiSTsBNZCeizMrP3YrzBPkYxHXKxrxD3+wvsCCtKJaF6klb7qJb2O/IZ+e2evQcz6OBWFYNW0/
hQYUesFI8UuEvRf1bTicQ/bN3HSmJvQ3WW/RPnepXkEN0nhSkCyAUkTXo0k8ddxncfYohVrXDEkx
8VyGdy17R0wOrEv3xEu0rX6hLIaQldDOW2g0X6M4vIgI9VPeGMpzs2yg6kCOIzrZ4OCy3+/FJLPI
qp8c24Q94cnOl6Q3oH0nA7cDs2Qh9Fpmxnf/Xm1GV7/qkvpga52iHrzguyaLBoa/5uIBP0Q4G6zC
L2NsPWqOO7S1ABuY4wILm7VfoauJ6NsSD5ZNM6j31edKt9ker6kRJtzT4I10XWMd7OPYp3/oiRwK
27jYhNkgDJIzOxEe0WV/q0tT+9ycah4hM/QRRN/IQz/CogLDAHExmCkRWufsVuZXlrS0fJoLHAgG
R3MB85KarFGsDT1rDGxfy+ydqT919pDO5HDLjJ7s3B5vJmXtgG0VOm0xv5NuXiJQGtPMerkp8xZA
wL34AH+WrTgViBvFu1oNo9Is3jiCu6L4VKXsnTdN9BURYBID5SDPMms5OVp4JJb6OXYRQSM3gw1d
0vSTSwIE8EpDQ5okxrh4mKNPzmqhZJf4jb1cM3eSPSPmL0qZMQcCfyPKJcWCz1f2kMKkNms8qxZq
e13ySqBHzB+/GI90MIadNrXfLQu3DJzrgrzKKDAG9n6b4JnpmsGcA5jEM/D4WfkraXNmR1xP2LBz
va2JzmHA5JC42RK5ckKM2LdXj9VKlxsCSvJ+p4971BcWvp4foVvwFfWvWYssEWKN2PXkv7oXHofM
x+Uhh59F0h9QQs8f1NH+tPUR0PoCS5xMmMTBMJjrDT5TglmptaAWxRsLjZa4zXHS6Oj9sAQIkrLJ
1GyWqRmutzC0AClA2zSPiz0jwKHcABJXd1tdimg6kNpYLyw4vAMIZ3lno+Tin8YmgggrAeq5VeM3
32pv+UkcaezwIEGQtLnI6ZM1VqOVdE97MH/njjFkg5bJnAFTn4nAoZMgxfhs9y8mrs1Ekf8RnVB8
qJmEcrogQyi1mnkK3Re3ZuM3IYZZm0TY7r1uAn2myxMHkT0baVe8CiJJQq22SI2lQyoxqN/jASw9
inZ7iQxvMnkrcTWDB8YSHGgi/25mLJEyrUlzJEsHwyD02sGP9E0vmPl/cz250+OzYYiug849qtcU
9Qgge5J60PIgnW20TNPyZxW91AtuJVvDjeqYPF6rCz6ERjSzXE/cOeZPnY4x3LyBA+vsCQnnmZeS
iSfdsbvgjr9gYILISgFxpAF1Vr8peHtM5itCrISLMheS2Jgz1OgWNTcTF8CIhLh5ZrKrw7npsKhq
JY5g3TxwJX7Tig04CrXl90dFRc7eAHR4Ph8fXNpTjEfk/tVAMupEgnauJVQTcCcUELSmf56FW1bg
G2jwMjkY/Xs1IT16fWWPDJjR5WYAatRVVMWeVC+Q0tY2+SY5ubLPQ1l8KJtUqfaQptFrwIAohQy0
j6x7aADCRFFY4xDfRezfTngwdC3sSzRWyTX8ooZ+NW2oPAZ3SJL83w2ILfTwdOXeMh/jKNSwWAPF
bQ08gjCNtiYSo/GMbh2mfF8P9MzRfYE3Mz9CRrZZyYIThctQwU0JYweH2g+zgJcYJqt3QMGo9Z57
WkIPr7FkgJSJot6BUStBHiixFdD9mqJYuxCyu6Ig9HN4lXMTELnDPMRaE9sNhZL86DZIXRk5kCRp
pQHsuQDZDmcEI6yAX5e4+xC09s5lEPxeGi2tkvPNFJOJPW7aZELu5gu+aoJTcoh9K0JJPZ/jt9iX
8fmmJWtmSeSpAQSnWn2omRcbq4/hI5c0G9ZWjmrUj1OEkLEBWEo+6jGFcc9UrmWErGDUBuV6GMSr
T2X6/LPnj+lIcG54XqFP79QfG45S+xQgcVxTCrSTvuukBsW2xOzQFR8Mm+QWz7KcnKchePNu7ykW
rjjydO6tXbhU18mkYrKRsG1pmB9K/po22UEfuU1Vzj8FhU1G6xHW+wClfNUnDkLxbFua7ijw+ytM
DFTVvJpXSKrFWPW+OsjnM6LjeDrpzlEPSoesGj3UQ3qTeO+5YuQ8J/kUhjv3OTwTf0Np7nEI0HD0
+p5bBKN8qUY6FGqFg9+FPTsqs2ZduVMktM6AkClMI5HFpwlz1Z05ghZjybVqCE2aZOqmTbpaZ+qn
Wy5aXAVsB1IJ1Sh5lmSCgPJYMPgGn/dpWWzmzOrnQgxp/RtKIG6Ol6/3/8kxhel6L35g1yq6Y8JV
e4287q+lZ+Yn57BmStA90dyA7twg88q6TjL3evNl1CvdoYoqDgVtFtef8Z3qaPneZuI4VGdCiy7R
+DvotNxb8AWo/zeDM+1F27W18VXbXbqNWMyXwTAf95upF123TjvvYmM28o53VxDEBqBLYJnDOrNK
AgrGBDhECa4qpCy8Zgay9NyX4NM+eD5TqGHd0rAudUzsvCFbJBRwd8nMLQgqVA8rvSktaJXHSTza
9dHy2nd1B3tf/G9qXRn0wmBC7tLhl3vbHEZELc53/gnvE8L0p9fDze0QWi07ZIrjUgFC7UxfmkKq
+ghJd/eWqGqSOD7Sb/kkpJ2aZdAIN1cUuyQL4k3I43K7muqKXL3/+ew794rsZi7r3bfAv9YzYCoL
VY66P0YxFA1cuh5h6iHK89yqXbPwwqxsTejZ4wsHVoP9u6SmCZ5Zz20TVD/aFH3Ol+jPJ+A2VCcd
T4cGEnaVBSs3rlj4HEI02Mc3KuGYqkTABVMHUGcESG/r5fsB6CsPRecsco+k/0dD0SFVGYq9DR8R
4lw/J1tIj5Y11EUhAfKkKj9ZtQ0MKPEt555Cp1EUVoU6C1nu6A3oNLihpiHboYH+6Ag3EV1Ho897
AC3nK/9O7TH7D2FI3fJKfpIQxMlto6GYwxJGhKYvJyFfyld6aBw39wQ9LSdIWWxGxu18c7abc/tU
gixZr2tskS3qnWsuUwlbzJalSSn7WqD5EO+aNTan9FDKyJ1hv2RA3D7MLl2i6Owq7o29tZDLgXMN
+IFDokFw4C3N0EfALypnaF5xHUqPX8g00o1CH1PUPv32Osnv3D5firkZEMk3Itp7pTReeeMtEpmg
4ehnqjCc+85RSKVsUYbhwlCppuzSI9nZZpDOVn89YO92E8rxx4n++N45wZluyBhS2Lw68hwj7Ron
s1ztyJsQ/GnZeiYDswGKS4CYP3lyujQ69Lif+x5JXdVyyJokfDXi8HMc6wZchsaRBJ4Y9ulbr7oN
UBohNcbWwuFFB87RfXzVuSKxfkhWJ1XEassG407MZKv+TesYaAd0R9w15WBviskj3fh4GDB5XCyr
wJTtQuCSbpZ60pBb151hXLyREL76ZF2v0Te/0ESjbMjPTcA2XlkDUYj9UszMsahnNYb5EENJRyoH
EpNE/FQiA2TnbIONUTMD39jEYSXPUpfHs/iK/ZoiGCQE/EQlVgygv+KoipazS4dnA1VVHFzIonTI
LHg4WE3/BK9wPwlp9qfra7vsa4r6JRSs0m/P55vTmfz9tZyGPPzeeEKh5JrbBznWznwH912vbrLK
7ixu0YmYyPyNp/ywHf5xt75rGqNruUEHq3Qi9JPI6snUPGfIO8RS6SsCKgTkwDFulRArqeU3UIaA
Z+8PYvSw+j1RGur2VdEvwULp3Gk1X9n+ZVJ0Qoam9Z92mhRJT0156022JFwh5qQ+Gz1upRud18ck
e4BFhadT36H78tiuDBcRiaD/81Nxo1GwbCSgTtiYS/eWrvOqeRJ1uuC8nt5+WExbfCioTQlYH1LR
LOrsuAXgf1YAuv4wqU4dEwmiJRgrbgCIPSKBh4u3uqyAMaIZLog+yFhEM0LolNa6tJZnq3mJG30Z
3+mTC8hz/iq2vcAal8Kg0l7PY6JFOR41UCJraUX/ErfCno0ehOrlKPeZ8TRFAZmBgI7tiazKoBhC
XRoLy2OoOdlM9E975TKCj0rXxpt83MVFJzi+C9jpguo/cAb4OWVy26MD23dEOGUcV7gFLJM1sDRz
XzCJ/6llhkY03DvhUHgt7DBJT/FLAC3Ul/v82cA9lK61Fs23wuZTKmgFuKtC7NqVKmvfabyJPtrE
Cb2kEZp2udQiWF+YTdbUKROI/B63tYYqzJb0DPFMORqUuKYIdtIVjprDDjMkZ8mh1BN7bY2ZO57y
z/PnujKIxxYjU3jL6KBPZy2hWPADAQUGQ723EIX8pnrvk26Nt7BW21j+aZQvgQAXs3BON3x+BThY
Zla050ov3rBxOCcRN66iY4yauC4Ux3fze7eb2yRMCnuGU+FTfTYpxtszGhnHnm3gM5tOK3hoDut3
Y1oRwztHA1KxVnVjPHarJXfYgAbf+leV0RcdBDZuZCAJ78XwVR0bXfCMlG4YQE+4Pg6WJJdEuL5/
nI29Gr4r1oWyr5v/pVBtPr4qwfrD06qTM3s+S1yYCPBK8imhcxIGfwYl9PsVRfNpKuHrEZp90p8h
lyf4C+HQTuByUteXijaNMCDgclnguECeRSIj/2WC245OEm5RbA+DGg869o1fsDI+a3NbPQ2ipXKU
KjYH9uXLLOUr0FPzeyqAdHx66/vyYHUr7gQ2BoPMSipUbTvMBRAfigwSQOXRdN+2pUgeMCFsXsf9
OSpI7NsIto1oWdG8LPExct0/4ChqqInKVoo/jWNz7jobsOiKvHREWjdGX7a60ZrN72XjcmDjjdk1
7NmNmj4r5qpmJevYNWyKIGJskP6GP4LoVhS+QlRvA8Q/tPZIEru8nYEktqMPZZzOdQJh2g9Ny1mT
slCyTD8sTsEaxac5Mp24zvmUmYqYmyWZQQxx+8uo49SaE07CKe3lADddvWH8qrIYWgeDZyaN29ga
q7T4IcS90a9l/cqhySYkaphD+xXEyrUItHnBWqeNaXXqTVfbzu94V/IinkFVoS9o/FBoatz/+UCy
ZfTIOZeKWg6SJhJ+M/v3VoH1U+ZWE1jzWv7TWZ3yfCjrN1ANzN+5N+sDD8ZSyBYonwWY/R7sP3OA
AxrauA4kkQRVGTyArux2XN1hh0BWZAMewDOD+pkW5+NB/ROj76KWdRbeBBOvk0gZ5iPvfRY3x52Z
VVG2J9/JGZ0YxLOi5HGsd9BH1UyIGlJWUbEi6ttZIh0Z1QVtHK/fYTzQwSdocztjpusFdaMo7IxM
3aOFP/6DGD6hVkot/TnJvGYllNZUoHdJ0aYLrFwwxeRMj6Kc7E9X//1FuozNsTcOGXRElRecaUs9
tRDyt08B2hg4Gpup9IZ+nUCFW4cbE05epB1LmKvdb18D5Ox6I3yP2MLbCMqK4JzTFirDj19rFwkh
nAxCO2wggNnAWZRHgyu9dVXR5bwL4l8coSwBFTudiUApAS30tkaSLTwJFNtFzNwfTpnhujV8vig9
WX1svZFMFkDx/288i34JuvoVpZIOWMPdltv1ntl43fVmLMCqHuyb42uN4EWQ2R+hUx5Z38rjIXOi
nyq9oiFQRS9XBuXfxNRC7SubU5NIeCWDl9/y2JTSbh3RPrPd6OmOaq+ysx0FyeaIPZ+fcndETyZh
8ddy9yCZp8M78iTgJZk0ZRlKc1km5AuvVHMVUwub98yeKwJdw5liFmtCQl2p3x0Qp3/a32Jw8N6p
C4dvg29NOcQls2m63prmMibIv6FLhVSmN1QaN22L/5HkTjDZkbaAFzQ0nNFyYwVJ7kubXYFQljnB
cxZjD9JCuIOYQp2VnT9KjtfLVUJqXjduq5AsVEtOSah6OWGhi5AWY7H87Uevmbj88LYiXS0KnHD/
HSD+NMuTzfSco4ee+l5oJXjZAF/Lriwgoy5Nq5DBdi5hmDoEUvHgMpRVDNgxviTFUlooiwP0w78D
O5NMxcpyZcilo5cQ1XHt6A8OM5B0aUCsKRRzmuN1/RBkhxbDUwp7xOWiGmn4NHV9Fa9Ky2odVi98
1aSttV92EDcpi5wipzxvLGsQw25UBNgbG2AS7FoBmYgJ3bDqJ25r9MLwFvk6z31XpD5jJIBlyzpF
tJ6f9L2wKnsL2MXTeb69EovXzF83avZK+LNenVCZat89vgeebPXejCdZeY1WbFfepKi/ZfE34sYR
+5CaSzbI8sx05wRuFmy38z4hR5BS7y2Qucki8hrSezP2eblQRPcmPQeo7TYHVvuEqTvT6btqZwiR
A1GFXRtcpyF2zdZzT6//Y17xGtxza/+gko0SI3KG5brQQ1wgAmsq8A/UUUG57rs/CvX2WPI5b5sh
Bw14Ee//q85EXoRRz8byIzOL3wuqpMRpx0iJ2DInbLbL4LxU8wfO+UzISu0PHYYU/JtPWJ6pXE8k
Jf+1yM4yn85X0hXdymPRtMbM/+61OA918Ek0nbBCvnRqJAlJP+WQbVxA55pqqUzVjJw6nwfZKEVP
cKbc5eumpe8eAgSPapXLIBwz8ynJ0UqGnNEC64EME+Og9t0AwzNh7rfvJYaFW+4TG87BEBtqQhdL
TChEm+eRs64S7cQgruW+MrOAhX9TcExl7Y85zl1ey+yBTbEHyqj09gwQft+56VHGF1RDSXETI0YO
f1zNKIDflYVDhrJaX7E8qrYL+M4TMuMKotq7labmo4VIlZIs4zb0j83F+z5T99Rltrl/yR3GJVJv
uFFMPX3ev/Rtc11rcdpOVAZ1f4cqnlQWs4pq+hngikUiSLUPb5TTmaUyv5CyMADI7x0A4+XHJZsl
JpEdZ2Nrrop4IfNAv4oG836qN6feywuwbOwy3+5OPTAayKKVzxcCAMjz4pNOmxer3xWUkGTkiQK1
PexMJrox0j/GFIe/pbk3GzQnatByFrAWvtsRzRnxrktP8IctJu9HZMG81Lr/JeXiFDIx7JZMmeRl
FGFSUnYqraJYafZpznrzeeUrYickc5ScS/ssp3nCFnPP/hRADgr4Zi7xCrKggwnZ8NZVl1EyeoNi
qtwUUS478/KudvL+Jp2CRsCPvNLnuZIFbZEIMHndqWZu4a0+Dk72uZq9Qlh3yVJ8n1iJZcia9pRg
NmgqL3ScAyq/4WjKrQG0bjNORRw78+L5H6NQ9JS8jE6iYX73dW2/G3JYFbF6jMV4COZ9E/STp4ij
LExXFu3OeWPCKPNM55lyGtbkIK4OmPdo8mzpImX6f+LwthL+pFmu/hbxThMnBeR9tvIgwms1lOhY
oQUf6LksJeTBVi14ONzkS4Qnwdbi0lCtUS6efmp7osjugDECeNsS63Qhloh6a7gbfmjCPs2KSmwQ
UhBa1wwVxVsL3caI/KmXxGDXxuf9XlNH2rEY5oUqZS705IC95/RTq9MJvH9uDfCOT57WOaacj+vP
/cX/HK0L/A0H+GRq/JePv9LJk+YFe1sudRYxZQAfiSKLsA0UMF1uclOxyFIf0PuIbVzocMi5AOAr
kj75WW9cXZnv3Me2VNMorIf6ZEMKDRgDTlJql//gA6spZJ0IAWbuivJokBTXd2F1ANv+LzXysh6x
/hawyJisXsElp7Hn36oUVxN3prBgMNBl5DNJaRVX9SU4zyWm0xtO2JyzP3VDrEiClQ5u8IJnTbks
vyW6CPDCtEQcp81ZavU68Bbhoo830bo63u34mWrpmMbzxoUIAS/MdJABmpfeF9TzJB7OIgqpAGMa
yHM36WpM89nvEdnYY7mHOj9n9QZNvT2ru8pvhSZaUnVAPz4Dn7Tm0lXJn2qyX4NPdqHLqdUkPKbN
7VvdXDlw+PGV3cYLFzP2SS8xIbQgMJ62mfBbPKE2km+EcF/6pLDbNGnMNe77i2lNc/cdOZVtHV8G
c56HrsSnCr5AI2l1ewX8I/CxzSC7QaLhzNzC+Z3KLquiVpExwPS8c3ZmnSYIC3QcR/o3eIWAYMXt
Z+z6VA4D2oL/y8nx5bTzWlRHgiqpI2KMLP/nMIfQ/wsfotBNqepYhaJrky1vKrVg+Knggg0XDTZl
S9eu0uiGF6/0FMwoMjnpffLyN8F2f/7p/k6QVol8dOqzvIo4ZfQGuqo+W1hFFx1/vgBa6/q6ttQo
eeI6AyRr9A+0k1srghM+hpo23ANHtNzC6qgewheKnEo1h9iWBPlFzQZduqkZTURW2geX+7iviEgG
bBpke1Co8123pRaoLjsPZpw2/A9AsGTWxZ98MlzEGeJwghXArxuVkQW1xCQXnCFMcfOQZaCS8DCL
r7q/PLV725t91xCorsR+jWiYwFzZMQHioHfH+gaBS54cOcFoDtZTuaTS79+Njth5AB7FZengXtb3
HrQwoLbnEZRdvOR9xjFzxDmKbhUtydkrx2w+mrvuHqSWwZLlA/q3bQ2R3LPYQk6zF654hP85yeTz
SGweeTHXL71E8oOSEIVXD5+5N2yOEx9d/TKAdvJ5wHoanmL3zcPVH0uxQDzGTizmqxWeyLbtHdZD
cfTQCIvJ7I8ClAGkh8X+tbzN+PvI3pU+ul9WeZRlYQztT5lP9CPOXuEIQC6eB8u2DPoBDrW9PGHW
GpO08JufKht4k+TQWEfb6u1ox6RSsmNTFH+LANbphBoW9UwPil4xo6jSnlj9hftY22rYhvaipdWy
BJenmM+snA8EXah6UZsNhY55mMqNqX6x2ULdOG5LEaXvvBGKbSGW3yp5uFZDUrdojamZxv8KZ0th
3GDdpje7mMkE2v68g0FnGl+rDT2T+kax8zQ+Sy+QucySL48DfK6MkfwjfYpxu5Sith5f6Eg8D88v
jyqzKUjvsEh1KCEVsgG0Lq3o++i3YvrSU6BIh5aVK0D2aNi1hlkiF2s9dXn3/APjSdUQIK64XBP9
cUvuGh6f7eAXt1ecB8GoieHCStj5NpPHv47/+w2+tYpELdJKrzGKz2IAUUf9y1evwVsz425MHoEV
pa3gPlRifpzbFUVKUyQQwZL02vC8FZ0gWYMtw8200vVgiGPkI4rR+xIWKYSL5kGT0+f1+v1bKRBF
zqFC7kycdWfbpAE2oA+OW0mIFd9ySPQQ823WAwa1xPyLMh3j/L8afaVpxDm2CzbJJjh9scalUtbn
QnAC/7Lu9aYvAw7TYjCbgPcZMCxAPXXl/kVpeBwZo6D4Mv512dbYBrfzA4cWUXMjU+Kf35L5O7az
S1ndK98h0+0G2AAdc4hMk4LC+++8GazTWhLbpbspUzkElZU2abMgyN7psHMCR4fKAg7padyJphXU
33ftVfy5jtNfRt3JzJ95XgcEkKJO+qvE8Ztu7bFf8Ey/IagIl775URAELho4WL7ioVJDGmqPuREd
i2zLRC8ts/jcudWB3f9p9EeT1v/nLxUXv0jjPp2qRlv5eLfGSrjZAlk9t2NHo9a4T6/bK3D5Wl3R
G4T06Vcm7sh7mFx8J1/jlFbDOxxtWF//BMv/AvadFWJ6NIONNvlEfC4F6A+KuGt0/HbN5rIBlCLj
YBExHLPnU1yMUvDsirVQEgEHnrtpKFmmWvtsHyarWEbqa5sqyHq/3ObbbulePo/ofC8fxmuUmoOO
ZM7XdilsIvVGmYQd+LdzJ7269Y7oyZCA3aAuUYrskY6r/XTtjoRIT86iRY/knM4I+e1neIPeDUJG
4oztDTOxWaRcXi45I9VErSmu/DBfhmfnjyWrxzDffNgLlB8eI6FNkzn2XVC4lb0Ep3r6ahYCJDjZ
7HQv/lDP/SEIk8Y6bgn3RKROJdjAmwRBRnPnSoPphY4mI5MDhk6kGJJI9wj8oEGk4bI9vPGTnlgu
g65r4UTGl35UGf64pf4AZToslXXpfO2/yUeB3D6+nMHtcAuhjsBkHatYnctT/aKy0GliXl7TonW0
wI6uRChV483qn8qoVuuJ7UEHHpc8fsJarwCMiPuBzLwRwD6fnt7WG8K7zDhpZs0ViUqKrb3Ewki4
GI4CB8t0+g60mfjmxVc19PJKUCqwVD7xbZCJlna4gOZtwjNYU8Wx1dKYzt6NcC/xIV7B+F2MO9m9
6DndFr9602PjIFBKJxPXnefT5HArPca1e2sw2E7d986OZljHoEVDhO6Xv5GZvHAX9+OdblFlOmnQ
qjpTv1iTq9JPXpC77cJGynD9LFjxgq6q6RBenCVusgn4t2UoYfPa4bvzWIleJ65Meuzw5PxY1vmT
mIgR3TG60A4l420as9TFHOc1Vi1pa1WwRHZSt0lnhXzwrqgZQkoMcFxeKwaKn8IJszPi8AOXJj8V
ziqeir12C9si2LjH/o131d4BktsuLCwJhpzi7pMH1OwgXmTrTnmjeddY8O68fFLMfkCCOBcvutzY
JRwQkupG+MTilsNdW1Q/g7Jeqe9ZJDy9fZxT//y6KgVLE4/04XnPApewvdCVZFpS0vOCN3AHhNbL
LNUqxqjQN8I8njm1bLQIBVHsrOz6fNsMgDUrmMYjiW6rLVT4G96Z6wxModgeO/WRwG/PPivejm/5
yOrl3c116XsHHrkaQhf5afykBLa4y5yH1yeoTgvhwB8cYmeoYues9DLROS5c5a1P8zh/d19LKr7E
YLNJkmNArpjyVm7vTBfrnqrPXdBpjPRxwsh30kcxiISvOknTmTGCOiDbuLgOxMvEmOHptrVzF8KB
UMRgU3vSzVKumZMQloZmi9TblithrjKJrEZgJ3xkOUSocB+jBqIlR+SYpS0OyprZl6e1mOyO9rXW
U+b078sQ136WbpIUVHrNH0ZujeI3oMf2fcr5b7iAUBH30KECvk76K2yxWs8BvdyWGvoJC0cdMK+3
ffK/+ahiaRf3paNXTR/mcqeKwc+AgZkgBUsPkCxtN5JMMNLUMwn9CVTW6thhcqlDnHrlbJaOYJnM
OTqMqdl6CIxNN9TgExEL9bUhB4rrUL4VtSKdjkMyWFBeRWLrzTwiLo/uSHcUFn5ZUvYRaNOSESjM
jXvPIll6EwQxMpS8u5ycTHTWQZNzX4qGY24zUxQnt9LGgGAXoh8FAmGwwrpSwI2cvV+9BoCW4/aA
hUK+eBN+ufzTbGU9SV7/A3pvCgTbl9vrBo5usJGm281uXlnFjb9spZuPlgks+tazmfmj8HkCsDzi
xeY0dT8FhkIc1BlMOYFi/5RzvumpRoLtkpzPt6Hyy41cx46+Gm0aXiEZ+O5WXNT18BpYP44YtGau
LhgtMSZTkB9UZD/VjIvPpIoDtLa8f5Vbt9SNwj3Y6xsvU58c3774xCmUJXJSHkjx7usOIzitEb67
rGr0ieU+xV7AmzzLkMWdeLiUGO7p4sxAdbZyFqO+mFARODtTMMejn5TpwTNwYsFk6kzFlZ2GAIDg
OMAaBIPCHEKsKSqaBgfgOu4w+ry8tajkkPUWJjBv9hziJsq2STsOGLam5cV0l6K/exJtVdMsUbS1
Zkb2UYUkphJJmSWfA8fBUUqELp8aGsIBpGJDXTghuJAY3nKNu2a4tyzjt+3VzifbJLUPvmbU428U
53EDmB7QTwyjn0wqIui11Dpc6d1ebacXKJvG3dVTM5z669ha2geY2/LkGI268z0WJYJJ4d9MXUXp
7tl5APlMCgf2eDjj5HeOJmAbtGbXJt7GMsFLJYOzz4b0zdbUppfsVV98puCsS6yYgH3BfU6unUaI
xBz3CU15f8FaXEO84NRuQHWjjP4C4Ag7cq7r0OGJuk14QWXNJnHpHbhPt1GyUWuGqeNFu3SmGumx
9+kIYVAtnH3xl8tCHMkrXmzzED84HPK+oipGrUqg+GB+Z61svo71m5o8MewMjjiZyzQzKOrgcoeA
lQrDG42/M6lYwhQL6DL5AUylZiwNqAd7MB12EIT5YMxk22KJ1qUEGrnWzZ+TWvfbsb3SXfTRHhId
Wi2CdujTN9fxiEDhhOjCZ4lvyih7s3xpTLaOdrGFVUEWPddb0PFmNp8D9TlgcgOECKQCYpb1iNqA
LMlpjuCD0KBLDjvv/ob+ixYNxoP1HuNx6ltTBY5XwZAEUgEGbgbfjQ+A+EcNiS39fNI/E9FKKxgl
9QNR9T6SOubQ/RFOe+ULq3ZGR+tpkWnpyeXdiZdM7iQGOqMHKnNEAWoLeZNrEkfZ7WP79NDKjQu/
Hxzpz8b8oe+3eWNpJIZsWud0c8kFfnlNVAN8RNIlod5xun8+1psG8DNtd4zN8/5UcM4I24AehRo3
Y5rU3teZvi9APRgiQgKIaeIFER536Fo1gKa7wlb62TB78WCkkY2DIeXY1uCTxa1Jx8wq7b6EJcY2
Gm0oDK3hBh2wjNUxqUvvohheI/nE9Ud5O7d4c+DlWhrzc4OD2fkW0yWKul8MEuKnrjoJckwuoDaE
Z615/aaM4KT6YOzQnJOK4EWeNhk/QAu/7u56o8/v36+OL6/MplG42r1eGd9eEPM/biJZ1SFV/gMj
IzLtB/J6nP1tIVPumNU7e6B8gcpvt+6qKxYpmCiFIsJDi69GZfuGLY8uXOyySQkwvqLcWIFWD8Ye
bqRQISe6I5qlkwk9SGDEFKx3khSiIqUbQePRI/EGCjUpOCwtZejmT/EUnte+APMY4svMjfTi89ZE
Kne3dM6SKM/4y+EzK0wQSajOt/lCQ0V8OL7TQK7TqWoiuPSgyC6kQz4AISO6O4ryacsq3xYWaH7s
WgdeotiSkfd4HlJdflmC8/RtBLKHCNaSOBeoWhe9OvPuvhtmo0A1Pe0ALFoLdBLR2pOF5/jRS+4O
RyIvy+52C01Sm0IzmlvEKIU7pOTC19snZyhwlw6wOZRUcJ8fmBVcJsu8/VbJ+v/hz+oQofjuwfTm
D6H97365z4IobL83e66jHAgcy86y7h7+GRIw4WQTyGft1kD26aDmR1UGCOiR7DD5vZzaCfLdegX2
jgFg0RBj2hRK96DCFiDVwbPR1CMmZ3veMpsqmyYZTG95h15n2BRNtkwetyEIDtw6bZZonb/D8YqK
wQG0V6KS+s7p+GLFuwU/G1LcFulQUVuDuFICdXcEtrZXa2CNbF7U7xPgpWG1CB1hd29+2iZKRJjh
BqVPTlAL2G65zAFvohyTv3CDOBuuaXt25taLOt5iW8ZmQ6zzYQNZ+ZVCxxmwHw9DB+ns49GeQmDs
sxW4BRDmv/Wl2bfBhu64Mcg7VF9QRhUFH1VQf3uyOLCM25yjSwx/H2fFIDfAMARiNT2+TvwPhlLV
GA+nYAQAUKCaklzk9nCr9Hpid9Zmmp7721wtIlsZtvFjQYB18LQG/J9Y9dp2g5NH6cDLesQ2IajF
i9YQVLDIDDjOlsr7rWdHwQLEQiPejOLzvqKxzK8qTY79eYe2YAsE9nATzMpy/PbTKargGsSXBOP3
zGx6exEBYOwyH0Y6x7pp50QjkD0MY9ZGWZWpgY/8e+NLsu308tdCBoyFFcEnOuWfk5XaBxzjSgCs
XEyAb+2vH9TkgvO2p9JTrlfJZZugsDyay0DVJV7GP+A7GQlm/Dw0zG2yAZZYAQEXBOz6xCp/MBjc
/IZL5MFrV8B3ul7WWssHL30GtwOuov1cxG80Y8dAW88WgM6IWS3UjCeNkt+VlWF+3RTOvTze8fIx
awY1ZFlzuqHpNNorCqeucJEC+Fq80Q4spq86H0PHoVsSu1+ZQQHzQtzwPgXYn/GuFOI3rAm24Us1
z7A/lICK8gGJBPhmqMs0qaqdYqZfcDNR2j4qy7spgB7pfg2/z2cKKjB9TerNozHuoJUkLdcLkcDd
Ima4EqJHdiysOwsHtHGnP6P4N/EpCsidp/2j3nJyO1PSGoS5dz68Dr2WRZhrtDdHiLShGJBK2Qnu
yfxQwohNMCWk+kkaIOFvAGfuvNKD3riKyZe0jI9zC+CW9qVc3yMCMX0CrbnnmYtvCr6O67AddYg5
nE3s4av8YkkJCl4TI6vEl611ZQczFYKkE0eA+VVZIkbP/ax4VLxkWkODsUhO/ZEqeuDImgWJtRwt
aXw2ySukupIWzZ/LXPVL6rmJDXHmZH16qFvWL/eaY4oajrbKSPzVEqTKUA1z9tXxD6Qo7QMyx9gx
MFcR32wYF90YKW67FSUvLn3PUFUJIqguSJS3nVRzCKGfsl9G6mqQU4+s8viYEgA9rDXDhzLoVzns
AgRfyQaT+M0nG3d4ZMxMNeth8bMJmp5USupNx9XDU2wBrXit10Bf8PQZcnVj4VA62XGnKvT0WjZE
IAeQbI1zwkmqWX0miqQpGXOI4csH0A2h8A3flo9NAqJKjDRvLnZSzRgD0dy2fQ5atM5A4p7oD8la
tVOvpnprcZsqRkkLKqdH5vWw0DJIKWZi8iPf9CMeEVjvJ7Tg4/E2oIChtou2AgW9yKCRCM3BGsLn
x6SlKVBD15/A/bIMRY8I9WUbXXwu514fBrwUElVhQtmP8Dv7gRhzdscK4BCE+D8FOnz7IuHgi/U2
fZuSS1rAPFaXiHpGpCSatdB2JtY72+Yg1ivLMDgELfCM/hbyOt1F3JcjFnX8flM5esBYFJvP5vnB
/q65qvTtb5PtmlbHlbfQnnDXTt52xjClKqU1vPljzgEDe9OJl3+8WIsDnOL6MfogbPalV2LRiHE7
n5ZbLRotrC2xxLf3xF4e6MrjesWGV0LtH5UuiytGu/skQanO+zTODSFGqr2sBsr0EjdRWgU2ywxp
ptcKwTMi8Zyp8zf1X00A6z/ePXm941mCl4ztW7enAkdc1xml+m35WO65aj2HuWTTOCz16U+ENls5
X85igA4kJ4/pQ+9JMX6hMFHkukYBwzJ+gJYLOhnc9EUV+5N5uzy5qLJN9TWcRIpHI8qzPvr/00dj
VgO4HF+jLbusVAvRiCEllncpALE+ttvmkohBUaDl3/8V+AvSPqpkAGS+XyFV892mOZbLBdTyKP0k
eCze0LOywDdOf9bDZzxQ/THqogA3cz+MAc/EzlgQwHx+uaDOFv/GO3qnotcB9E2pRkAEuGWkMkEK
zaH7if9sWmzIyje5lK/QAkZrhGn7/ZxXel2mQM+gJhOl9vp+XILoEqxChUzt14Vad+7ENuyAnVB9
mcUOi07Fkn11y47c5IBlcn9Y7Q9KF7OJMS/Xooip/fdu++izAED5a3z3mbGY3CiX+ASOTOy22Dfh
WPMLD2ya/3+ByEMQhYk1hG6QcNsAcOYeZL9sGZZD3m+u3hDmrClMu86p8YespMW3Qj7zx8kxkin0
kMoNnH3G5hBRRIgkvWWvVbeccZYD5KjCoeQJIfXdBz/inhQjpEm06shWVzgC725DxvKiotxFRUHp
GL5IQUIj7UHjIfAeQfUoJEn/Bv4uyVvNjxRA0hG+Zsyx6jCSTObaFLLL/Okru1ybhhRCSwOq0uyP
1qNXGydS7/HMQPJA+MoRif2kj0ofDqfAQplu0S519Z0WESK95NbiafsAyA0uiDHadVJmFwwvM7uA
2afMG/O4pvFAYpRb6o1/j+I5/FcCGfA2LjnuODtnTvfenFvE11gcvZJry6OW/C1X3SS4Hz5ltgo3
282p8HXZyy53k7W8Mi0n4ATYY0bhQkHaBBhdXBKOSD198070IILm5NAxnuPyCXOuME+3ApwLTKPT
sCNiIz2h5d1yWM9H64qZiDg9pHFc48w+Fp/2vnyMGuC9f8duCjIG2aHGAwQoNQt28GYhgPxUR2NK
cwyPFXK05FICQDEwiNBoIjQ2LaqaW+nkNzdeIZQDHWHDHSWz7hABNnLQ6WgylT5su1lr8CjeC8Pt
5OoW6+25V4Y/fooZuh7vXhEOhUEsihKbeGL+0WwtWA7dwP+r/Hn3UpNs/w9ka2/EKxM8DM9U/rlL
u4mXcl9YoqGgvHJUlRF1FFlpsxwZmidpaI+yJQQ3wigLCKhXz1fvOVUcIICG9tLIXj0jtNqU8Mao
IBr5s8lJFVzlW5tHIzdRhvbr8RAoqlr/+N5DWfZCeGm/c7X1CCfzHSR+fapWOFC1RMkK2YC4oFNp
AvLT8bACDjeMGYooiAKbn96ubTaHWEwZUkYd/2yp0ZSngi7LK+66m/RL7IzamUnXLGT+a8GFNsxS
AkbWj0N5yhTO/qQjz3Ubyxg2hbm53JCVYxC2x90UA6rLE20reukR3fr9JVoDQFeBEkcZQZrT0BA7
9sukERxYFjyJ5K1P5tVIfhcI+DP8F61xgUCIJfwLR3xL7YTWCG//cQgkMSZtjdyHS9sjpO8ceoiC
LKB9MUxsqp8BZ+wPQFtdJuUo869cXppaeH9FOkrx3+ROmIDRQGYgLpDduA1KspgaXaxL81OvQ0s8
vRJ5swp+6Rtsm40qQysxe4ZXi6u4g5L/rhpDN8yCdkdO8JLhZNLtYVq7nxVLyhLbNhqncA0E/Zp+
9zXOR/bXoDRcUnJt1reuhZsZ62swT/UtY7/1Q/6a3TQCu50SSYVu2JT5WM0X/XdqfofmeBkrzQ3r
4nXb3mhiNlBzp+Sdzlr1vzA0cfdOogwJjpdfLdDzqh+sgypgWgmRq2S607lzInPK13PHjjxrgcKz
d2XhGfXoieqgZZO5nMk068Lgfrjoiv0aMKnKtJmD6Q0YjNTqhN+JsutxndAjEmVcfVyMBaVPrqtQ
kmNkHydBPH8zySRDF5RWraNOw+urK2Y/O3nDK1TK8QfLv50qq5zX9mcFGzKjTHh0XE0vXKOnG2vP
stwhedZmOHbPDIJxPGU5QqZLeG6C1hPQMEsOJxMUHyhF/BT5nFdzCELrOuoTqEYsJNC+xaPIr5YR
w5Ubf2q8oiqgIIqHvlh2S0DRRXp9XGoIESn4FIzxrS0B6zXo3A2TSowQGiMrhQV2HlYDrDS94G7K
0GpgwEgWMCmx072oy7knmVyTtkpqaF37x+nwtxt+HAZ04KUbwUQzC0WAtOsFZw+d/21REyhOjoq4
cwQjOM7Xf5JeLZpGt4FyxfCPIqRQDlRE8XRPPTvqZ+v+wpBDbo3ANMS9Bn61JaU1UJs9v0zMymJK
aOfx6NN+d89P+v4Egt+Aj6Xx0yPyBM5sumOf1DKV9ASXvIDHYBeS4e//UHJ3M2PKA/xQjWwvYukV
Gp05hIXttf4F2rBuZC3iivXiFL1TttiUa8YR6tCqSxBPuZpMcPMUKTKgKIKVXfWM36niSjDNUdGY
O4pzkVHIg7+xB7sq32RpTZTcfC9lTiVFx1tWHDUsPtei5yfN37FKf0zzj2viu1ModLGA21aECXGD
7siF3446o8aPRGsCa6DQiQDkQ+RmpN9vzNWhZYFsvj751HzGv+P8NNMMJeKBImV0U4ose7uesCJF
BCpwbR5RpJCb7yO0xNKMvXkmFtyhnieCCEB7pfyxazpHSd+1Lhk2D8iYDOQZLOOqw1JRP7ytr3jw
kd/SF6jqSaXErztzeyOysL9FPVVR1brPcN5c/4Q/GBVHcnH7s/65rXwj3plbqbiOMEVbbCOwLB8X
QN9BDwIqi0AXM8LUKeuRaCyW9aDytF3WVFBrHeybI4yn5/xZp0Iy1DaBAoWQFY+kLmkTw4AFCHUu
pMCRq+cUnz1v7O9eaDmeETIU2ypabL1DMEAeAuyOsBkgCa6shqwfr9CLYX6GfuM+2sKjJB68aqX3
V6QBB3ZtA4K/UyDTZ9gihWMyvwhZdWaT3gWeqjYx1VXQFUa9/uHZg0JBlbjemgQ0BXxXDwU4GATI
qNRAmEVYahhV1R3s9ikm3Sf45J/w5Mk1xfWvkz55xj9oSlWyFQePmGxdck6Ysc/EkD2DFAg6HcYb
FWlTsLpI8pvUIOPmMbNmaijudNJb/2tAQicigVrepU5IRLWFe7afV8NbNrYkTCkFfase/YpVfJmr
rcEbfoPDGS9vQKF4STalibIgHA95wvVJ+B86HqRNDIl2Ul4XlGwhINQW3Wlqd12Rcq+ilPxQYu8K
AYX4WnBeUMVh0lvzkIzh7uxRmzgIU5EwV1FtyuOfv0+UfyNofY4aYG9J+n5yC8O6MXYzhsYT4pdm
AFyySikn6+xq7y1Iznz8zCtAzq2tFKiDinFwwjNdcbvu/i2NtPUMcBOSFzpTBlfpRNYuA18QDEhx
em7FsSyVrO4VU9/YR2A3JSzlGdT+lTbCRfvoKDvtnIZCbwZhsvDSmzVpdj/f9MaeUKjVc0KhnNwW
Gv6CE1mWQ37DTEmZ8x4g5/iQiO3W7fCIvf+o95+4YukO+Uj8LKsFP1YPKL7yvsetuOzTOYTs8AXE
guDZqR1+F1oFpwraCPzMg9HfkZzYB/tHubBXv1Kt46x70BCAy85vUOOJGOrxYn8ayyTPPew06ExT
9bVWNwrr/I492Ha3k2rufOiXb5rc2S4scwP2hhbYX3g4GS4owN2o5gELOF9TWsgTMu494ZLk73tW
P8FclZjpd6I2gaaYlsPcDlLe0skR5LyrNGbLejDFDNm4R160xr9RofAEcg+37eg78O3wsVRXHZ8W
r040fYby03tnk0H0v9c1vKPhhzX2fuRbjyBywej5K+bq9E3rzhNAsNbMboz7zQyXf9KPsNZzEEn8
KprrOymZK1Rfiq6w252WVGRBSfZzgTprutuGb2uEKvMm1c4wLefNoCLIjaF5qhJwggczCO32yvDE
9SG4DPZDkYJiPEiCRRED2xZDyFHYnratRevhB259CkBGH3TP/LkVbouY/s4vg75IebaXarWYPmoh
dVcoR2MviXxpy2MzypUyO0REqeZTHpgy4eHPrCxYduQ+lEF6fP3Ma0P9ucXjzIN3NvdV6inzINJ9
2gpZkfDrq+HgkOlYDyXeAb2DbWpda7kRQVkpYmgGq7uXUw+sKpuXgXVMydgP7BvPBfL/fbPdD4ih
/Zp4f8/Z79ltPfYm2Z7jaKTpO7ex5f0ccfoUGK6QpBb+OI4RNfRSZC6rI5nzz+P6DHIX+Q7nSJFW
Gv927ZGhgbpuEg5FButht1Q1uAfvWMs3pNcdgX2PNP105uO4CDnhge3rhPnPC27vD9KunICh/kCf
vPd9h0O6GP86TT7NcW2L4WfpVDXZdOEkw8mIGu735bi5g2r6wMWwHEELtZmBrjTRDWi779Kn8BrL
ioBt5GPmF+WM2SY3QTlIWmMIgpHdlA7d3tvj+pNQlLqWRHtdyr/QmQssNwuaGvqatsK0HxOZnMzn
hf36NQ/x+DSMHqW366dl4CV5DlzX3QgLndZyY3iIUEkk4gYYvU++YhDniOURUH3Nw+DdRL5a3CDE
OReQ2Fw20NUTdv1t0mm3khrhJzuKsiGmMgQBAH2iWV7kPge/qYv0nACoUH0MWawPwduWHs7wJubl
ufECqSti/7CBP4VcaPcGyaNvB9bfgWocf4mflYctcJbFNuxNt7JaDNeb06T1XUWg6x3+JiDFMGLe
1iby0kDy//KvRk7jprz277nXoQWPl72aVnBVQTqYRhsA6A/5x/Sh6M1fWPLsMMjvNwSyhOQ86lC6
UmlOOEJUhKtqVYCIdYFkUANig7jBXK0DlieGVBJr7VhHvmJupe3NskqgbJ1GtVBgsdibHNK4ltuB
mqBTbjo9AZiTqDiz2tzIMuBKTzGQkDXyROjwle4LjFw1uBz3qcVpNDder1qiSbTDkbQxmd/JUYJx
HNuepakDZe2KoNAouR9kcgnfD+dwlzSZ3RXm5SXt6U+rgBwtDIrBPtRcTffelQRH3YBFijKEpAqz
0ccrtTRD7gHI9GpN5FcL8zEXRUj0c5l8jZT4WI8mWPfg9Pf0T72YhKgB95GHZBDa51tIaqWSQaIx
jfWOhQ/597+kRHsHZV+zc/NFsdmHByORY26zhbdMX4lu/Hf9EsBPA5+ZAXyYbXy4CM/qiA5imbHb
lOT96EDMazezbKycP1W6Bh2LhMoPqptYtSRSpP2nZmhrGNn3GIQJLElqQE873UITxZKeZl+ahXUa
Bp2zhtWHKrpFBaM2fKwas55dMkyKyML0hkyKd7Uk2mGwRI1Hrs/RP4VGMD4Zmvlc2V0dHGakWeR5
iOkvqQ0YNsY3ZKaBIWUzQYaasc+bQm7hxd4DAQ5aNtO//89D9uT9HYirttUTHlzFysD5lTeAVFrd
uQ/J8+d4HArrCblI8oefyx8KPF/3HwYsd6qe5VrTSCwm9T9i8qVTgmaIrIKKY4L+fSWBt2FjXuY7
d8Ey5sq0ImAG34Bby23cjZIAP7JU4+h93O6n+Id/T4oH0lx7Uf9bvGUX0rxFkd7gRjn1wXjZcqgA
p3J87EUleyy+U4eQrQBgOlNEzu8dpzFWCwiYx4+PK1V9f0hKYb/X9JNTtyjH1+KVC6fGiwDvGctc
dIo2FSF2iiorZPYYIPaMdRG+y/LQ8HzbmthggXLWX2b7JEdd0ARNEzov/QkbGctkMfXiyJ9IUHMX
+lUx9DrSQQ08FC/cf8uNKhFVwl5T8hjxgMXrr6nnr4aUy6tgvcjCym9RoxqpOY4lPmhCVD5EAeqn
QIczjF+of6G9rrNdpLzIaZfV3HEcwZoQPF+HFuzTFyH8gBel3B2TPW+C8n/LUM+MfWiVqh9zppW0
inl5WdIXfM3f8tkP+zYWCfqeebKTDwn/dF/7M/tpqqec8pS+xEhbUu7fbCjNrk26S5mcCcfC8n+M
rqUpCPdxPH6nAh36JvB3MN6vU2eallW2hrFjLmbST1PMG2Tu+iq4hR4Alxm5HFeuWfCKW60B+WW1
49vZTerFffijeuYBaW1cTgr2474KcJXARBAZTEqvNxX0qDWroA0P4+RdZ81NXxw+Bakz4quS5a6e
2DfY2++27V9+JE+8bx0dzkTZarAJqiUN8lSJHoeBI5JBvGyTt8AOQvu/IThuI0o2SHzjfA1L/0X/
n+nUiDqzCZg3PE4X9hmAxDUkUaV6KRgomsq9WdrHNVzBb5+oGnndcAeV/8s9DK8Efx7biXbjFiA8
TdK4GTjVFz/oxVf3AL3PxmGN8eW5M8Ap2iCUCNzphKszAZYqFsScy6+KKKs8a2K5e862DCAWURAX
Jn/Ci7YbA+7Gg+OrXe3X4bMGezn6Wt4Reehs5YTSFxxxbQ8eRRmvZwJ85zqgH79m31Y0azH5Fje6
yZH9Vc3++dEXK089zfCZIeEEBs1Gral/x/MK+XS8G9mPqK9pxbmtAxcfybsDuKvyMxw4uc89tPc0
EzGyw+oizyHmzSvA3RBqwN+kJKy7RSFeYTcRZ7USqgJUIfP/8jA44lE+RwQ14VJOx96V8KAciW6+
1R9lj9Iq1hw+YW9MXEUTulswYAJj6m2RsXqfMVowgJtuRdHurbe1VdXAABGjcPjUQuSYasYVokCp
8L9AIvbhwDfwXh4zq/e03zNDfbwNy1I770tLx5kxSjQJ+iKzk4/iArUQWM5Vz2ljc/uI1QIU1q6z
VLcJ2DgZvdxfkrqjcw9NTzWuTNVtlN2r1JiIoKogkqfyUB30Ue1yHQyrVTorwA/Lf86t40A5WQYn
IoHfkdbvWbo0Ip6BvwUXxELYG19oAbEoPf14oPRxCVFWSqbJfMnWPMMQQS2/aj/om/lHpA+7xHaD
+7aphFshdhPmOQc11zDbqgxxherJuJtp/bv9n+1T5orvHjvo0eKU5+QNBtSsUrWC6LUaEuoujhBN
UMlizqms/08J1AEVRlTAQsrHcfIFtq5eT0dl/1W/JGshGOYz0HV/pSNmYWV/aMlS30Jb//LYbK1W
MCvufT92kTeCuyo9s7kGK4/sLphiFMxStmZCtBObqcyz3QFc7c4RzA8JdNyU+8Sw1nD7Qf7ziMTc
jtpWllxoSBHOugsQwdY8G17iFhqEFQO+vzTFS/o8b9sBTLWpTHEzCsRQ/D1GHcvJeWnE2ceT/2gb
pKptj8Yl5b8d+zhbXDOuqDNZfuWk1bN8+/rEHxuvXfaA9bcc6Mf1VDm4wVf0H9LiB33C+xCLYsIA
QBVk1DrVK1ORvXeYShXEPDTsiKW32j/xlmft1JEcSNJvVdG77WwetuJhBIyy9uCcLhujvXKGqmjm
I45WRGFmw+WDYx7xnF7aNhSgfag37iGubQlqYXed5oxIIQd/weInrmBoxoWz0RJVZZuncnaUc429
p64Hdsbf3Yb1OJ6+gvZVrx0kDhXI4tP8WDe1kvxuKOjsGsB2tQwRjmsjFN8v9veXiWOUhYwOdh2r
f8aOWWGPglCvNkgrFon/xR4a4594E3dIqKh1EAWRwKfDEzuUrah8M24WpuSfZNmDET0vfJaMu5lY
Ai9uEA8xxSOvs1YroyN68h2tc4H6lLrA6hQsgp5h8ShDldUvPlamYy4j4X0FuByaYYQDn/PZ6B0+
haMzsgsiIucSHeiA0IiF8ACz9rRcYWHSZf1YLfsrDXmxoTgbwcUkbtU0E9KTN18iGMqWpMAQSo+a
Dyd9JezLwZXD045cx5a0xOrb5lz+a46zH1R0RI4EDk2hopyFpRazgze80F+nMqKwWXPMWizKUdVC
yXL6vruUXdcp7uZSAroenSmqVROLJJjJQyhsoSarTTSgEM3qoOrShuaXwtYZpmkwbga9S4iAucds
x6yW8wYYWDJpRxacVnj1Fc1T0u2nRgThsAZhtDkHAkmJfDnJWb9NGUFbsL93XTJNYk2uE4izKEYp
ET3zLRuMvUlOpNlcn5g/GEzPkjxlADwVV1RJEwVg2TjmKkWcG7SVrHnvEKzzx8L3/abc2L9Pa6Bv
YtZ59a281t04qFwNTO+1yzQEvd3CsZt1QmiWnGpzV91cbpMRo/xG0bazebY7qSzPpH3XvrJPPFbN
jSkVKN7oKvsJLKa7LPFHvPYEGtlegbK4WtEIyv5gh41HluqA10v/6S1ZFpIDlC9reKe2/Iojv8HU
9pVgyMhA1jxFLf9o36kRzb5yTWNidNlfprbCaLzMF3jNE9Fm1yha9ticeqXd19wv1Vh+6hYFosH2
9ucyFNyq7BqspU7pN4gJni7XcioLpW/EGNemhiNdX24BWJ07ree/IR/fEFFy54TftexAhXA/TwrE
5FG3czn5nvoSsS1G7KjRTkrhHQNiWaCJWlnVs87bI4fa9JySVtqkHPur7Uu22NtVGtapXZkfs8Ha
QJ0xGY+hQFIuBUTkXz2LwI3JW+4hZtCvqrz7PH33ZqXMIekIwgwjw2DoM/gY9K43iLjl5LzMeEHK
cJsaw7gV+4NLIKCYc2LAx7zsgAqu5CnR6XLjA5sKz1IY7O8aHut1wxW0AWU8NaSgk5ztKBux5UCD
HpiDGTj9sEeM9fSXRNmSoH2TwQqoRdPrF++SIaC7n3TXTYyRzqpnhstUBGKri638R+wCVZW7Smfw
VZQtG2anLWFj3+DA4vdOhBWeSoqglE9RpFuVDAXzOrN/e+oqFgc/a85KU6BQdOhfPBQKbESKO1xu
lvjW1Wb1UwiFgT+TvZ/j80nXcl4Z9s5APjiKmNuy2L63DNl0RHjpgitDpiJ8Vo2xHL8oBkCz3dkn
GXRnNqR8ok0ADYdr20dXXB+mbSmS9xsNHrsEwjqk1K8zqS1WQh42bwmTnRT18Ub0VDwMwAFmRxku
mIMnj49vn2j5K0VfDvLpX/4kMysmEzcQncEZOE8mCg3BLbmWeFVVuHP6Y7OukEByEXa81Q1czkFX
ysbeQ4Rw9v2yiCTtTrefZOIZ6CSR4RJAgZy6CDc4+5s6USEye1919HDLeVbYvMMQlnGigFQXKHbn
RwnaVidI45Gt3Jrs+iFR4Juk+5fG/7F1RrK+NuiUdHqxr5Qf6biMCeRtl7KOjmapiR7brbQAELUk
SAcUcTkWjmteKy8dQ2i40rcp4nCPe8xV4CbWFuZygxu9yHSv4bf1XIf/BSbYPVuXavJ+O8jExDwZ
gII5j037phq9MSIkplEFT2XRzCU8u8nxQc1uKmgdWB9nztc6+ngM2E6xnFJ3FCPAz5c5d50uEMO4
czWCg/7zNltxdfBYSiY5SJunigUibgC4zs6CUZ1b3QKhjFPDTClnVorrD0jJvdDXe97xy7dTOBTv
Zlex9BXwhW3OhvDSl31gb4oIrRTJpcVceNrb7mOmrF0qRApzaXrtEy8+4c6SPRdMS37i62A/dgER
rpZL5vu6pbN96JIM6VHjrES1Zs3r45YimIiWC/bUZetTY3f6S1t6hJjZPlPNAU0oDVzNXZSkKTWZ
ud4mdfBUjpI9IIM20BgDHSf3jXJOrL9l8GIUdjBt7q9LGTmelqJ/ymNSeDCYY0V6SYjZEHjDfcTk
DnT1Z0jF3cYhIm263akQS6+xYnERytkv4iHyGBg4pd1e5rdj2Z0e47h2HjWVYBTKJqswhmm233fm
NV1fp0Q6vpVvOHn2v8JY6pARWX0DBMs2FIgnc7KBd1jkVZHfgcerDTnYE75D9Bq7iKw1d9i83cdy
nRfmKXhXUo05IvQTb9riHRj1MauLJHK+kbyHX67L4GWMnE83vOmXLJCKO5NNaOAdddVOcNFccJJ6
8WB2j09Z7N/cwF15BHA1mD3vkrETEP6LFbosERlp/xwHfhsxunlJUpoyhsMQ2ZTEh1r86biWzuG4
DcJaJrc5FTzeox48fSMsbprMggRrFT/sRyElG8wsUYIalW2F+H8TRhkePLC7ikqppnlKJdN617tc
nYcEr2boWNkduUzulY765ftYfVskMB3E+7Pzuv3pgFhh/Zg7XLBuSQ6dJGOKRNjPL0eONTnwp8ob
2fjkR5JH6lACbIM8fTZ7XQECC+bGhWG5dhLxlgRXdalNBhIgkLud+VipIzKDu/AdodI0DzV3DrfP
CvzX2DfNtGJ785z/+Lc/CMyHrn7jsGzmrySq1Ivv59XMG25O+3n48JBcPU6+asGWf7viyovgT14A
BQlctp1yYkugDM+tr19YCCohqRAYtKxTT2Oppf5wilujKQYbELOx6FeEpZjNueXEC2uA/GbJ9m1P
Xf59SSVkyOde14ovxEAJ5vcZpyu1+1zyOjsznH/FgQdWwvpDi1M7t0t3wS7VO0QJNF9a0YsUBPjy
Kridgjl0V7wsZEsp9A8JhzYwL1qqEckGY9n7BTNe/AKOSfz566FovECFMbI1ZPa/lTxmi0wCu8Qk
5tbXO43FPHKgIvdUp8BiHYZU30PR0kFy7Js4eqNP+ZWU7afy/ZpgT8ub8DXf6njo0rSpsx8z2c5P
B8G/cYym/X3uSt0gDI7AXtQ4qhd06vmCU3E81+q4oHHrGjzk5QVAkE1KSLLDBxDtdtCskJew2YY3
/8wY/zk4ubWL+v6Crccbu0HlAO7nXbCSgueHNXhMYy0kpzq1zsT+pNBgaLnyAqY+R3Y4ie97laN1
o4eI2CRuXA5zDbatk31p6T380XxATxB8sD0Vgb88I9aHUlCzpenTsTUTvit2+XgEyIb9/GpxDNwf
oveZtU4QzWBc42n5PuRrs7RHSEPRExlUpobgubBE/ZI22lpy/JQsDQZXIRTBSfgupVAEvsNfWn7G
F0z+yWrZ0uRlqEIt+J1K/rTtiIoLBANG4bZ9GbhSQaeTk0wY0GF1shzAHd4p3JVyAC3fEQYQzQdT
jh/KjxEw4Tc4Bj9OeDUEeKJoJrCj1Bji4qDW05+MIszjvR8b2fM5LCq1OGJUuWNsjpobcOtZUWgY
4hTHZIZ0LMckWa/4gJl1ToFNdg4ZTv8qRF/ZvpQDk1cLlibwgbepcaABJxs+P1M4y4SoXBjxtNSt
Q1zJZSIYsrKlXrpMYNL4aV0ppX2QpO2Jro/M7oOjx5LMdg49qWlbt7yVg8svilPSpL2wU2JNL1Zl
u8ICBberjaU9jjC/4my7lWwYzadr7bnPRyHrEIWrTpN7efi/2aOY7dcYqE89v3jVUThOLl79R7/1
Pr3n1xgRdQelQTBs47RMGpMlVsD+R3FlfI9Qsc+fZK3wufIgx9Ir2RzbWj4gyYV0dMqJ7PueEb9L
m2zaUQJiziB3gT3RdgTXGTqxaky7l1DBMBg+lKxlHvfR3JRHdV6uuwT/JQQw48SasqPIt39o0p7o
+3QViZkEoHsI42jMWzeJSqnYxRMALlQYANbmpfcB/cakq5OrsXiT5XnK0IW4SkMtE4AIzT5D61B5
/wDdh31fRhFqcyGIyGfaUCMgudvWmbOI3SfXxtRutUZNS2QXU9XBzvhE64+UHm6lGAFN4Nc1TcUU
J+JJ0Pcdk8ZPVoSzf8KRcYc3ru650Z6dI9xeIGQvUZmsgc5Z2GRHw6fQsA/8+fkV6vllYte2U3Vh
0lWgbiYON2/bLh37j53ztcnpokGbzv8d57s+gsG17hzxGFXFuk/15GlxNYPXBt4TGr8sYcEvxOp1
DBuv+Xb2xKBedDWYI3/K6SGk6dceEBaNmpIyh4ODbfhxF/hJqtVbAj8RGANP8hNcHIqCWf7Tu0y/
btsdwRgudriwfj3Bdy1f7JW7ETLwMKOFWJnrWEGF4vEWTXkVVO72hcFg3m9D3J4gngUvAGgMGCXA
szArgq2EWKJ1i/uUg81GIps8eFx8PWgobZ2VEkp6qj87zHItvqw+4M5fMynB9W2tcoppcODhxQpi
/UoiaNFMgbDs/Wi+F9KVyZMtv0ciWlCAKtl12DB8/U4/W7C+PHi4bsQCmNBPiFo+nl1sQnEBaWtG
sWDQiCnunelSH0A/AiYQAN1kdmTNmveT5zWOYlUnAljYYidNj9R5tsrGSzhC4w7EvUvDv6nMbO7F
5UUh1I4kUQehv+IBAVZLf2ojt2DRE8dYxNbaqU4XpPZrxQK0Y0srJww0OR7xtehpzneAON2pnWtv
DbcIDi0BTnRKWZlyZNs4h1F0z3CONolvGd4xm0VcdqAp/ljmHLo2TET6lWdAYJY5mH+lzF2u2ZoG
K+cc0ELei9tvrpJbD6kRzxjnLojer4REwT6gyyB0PRvVdGICImbiLi4VUostQE0aOmj4qlQN2xJo
b3Ejxzzr8GPkV27uwEeKpz9GE2Fl2uir0KfzqZHI2Er2mwtEQRRtvboHBVzqJhQBIHgLXDaal7tr
cjtwJW+hSyvcyQ2EUpBVMxlHlaOKgtJODaoG0qCiqXMakf6YHpqyeXf1t6waS/lyMXRPsTYSGIy5
4ivA/+kTXShnK2gvPGd0dHnunUIxFgt2RIWudNDqaDaXrKLFu2JsWNAuSa9srZ1pccTqYYEloT8k
xV3GzOEedGFCBYzK/+0MyYtKk2QVb2JFSl2eQqgG8xMUcAHin0eJdqVzZ7QDLKvtA+RBqpvkBdfA
FRC17PvS/M38jLYusujtdLmiM6GzM8qAjl54zoqFmbA55BeMIAJY8rFkjNlm+L7huXut2iBBZo1A
kC4K38uiVKBZYSQ1xm1FRNo8yQexM4nwOGvS5kSkMdk1Je0jXWz6QZioRYrlR/BgZeulljJ8O8r2
TCGG8CDidHtoG1ukpdexuxDbpQLhR0X8vHnf1bw3LkOHzYlON0ilMwVBZCqWc+tAtNxKMOIY6jPa
Tr6DvlHtPHrLXfy3sDAT9uolbJrtUYgJxRCAy0+KCS//b3RRP2amorQkO+cz8QegWyDLqjud+/jK
0aJd/vbKiLdA+/P8YREp5G076TZbtUxunPxLdsadOtwN+cU6Zhzn28iVd8XWXOvyQKrdEe0Si5og
jxXoUzNs20pxaQAoMbowlf34KDbC9lNKwTxTkq4m1BPqaTsr6Y+5zvOarmZFz7GF2iYHwx5O9MRY
NwfqetyyZkjGRCn968tvwypktTcLupIoCe00AKTonIWNqf+6cu4+OACjzSGCdI9PGEDWziuDrVv6
kx+71fgLn3YdLYox0OECCRypRUaR8UuQCdnNMZIWBQQ8maXYoZmFYAWWgVu448vOiN9bUtYp8hRR
yLCoSYGh51hZ7R/45RWD8G/wVTBecYXDjre0UNz/ZnvxfQGcN1ivwmkpEhXUP1Byk9ewullBYn0s
2BrA+mtaPtD90P1ozo/6dKJpAjIv6oCNi+Rw6JA2ly514kZ81JwJW8hZVHXpMdxrMJVk7E5shq42
wa/8av+rOcvqmNcv5h+NJwdfvVHNwWwijTZRgQ7HCKLwnvruNep1CI4aBkNc+Svc6hez7aAmNS50
oJUZggcsWay062SxMqUcjOCeewAz9qNwePvRqGluBQSddYSPzuLIS+3OCGPD/1iVBX7c6sU5E7i+
2wrPxkans3bWfm/TTg6JBzZrg8o1MmE8zY+s4VLCJZWmZLUI9jexOVfLVJGW5BiYthvBtokRqnch
sBUO5YNGFz0XyK2FojxXsfmOB90nxS2IR2ansypasqRjS49akvEbDPmLbHJIMKaFmOQ7Yw9mPZ/E
ybQ7xdNUjqQpUU8M0j8W7qt4fDgKIQh9OWtaI+PpNmESTrY9WjYWEwez8moy/DEC5KFU9XAK/SOQ
cteTOo6sV6+HQQARAS/CnC4j5NSLL9rve+V7/fR2WWJjks0X3zjPpBJXWBiPwY/1lKq9H44khIc1
QTgDGHut95d0TdOAJ25LvKreWgGxRUuX/gjsydkmRkqPY46oLJukE4GHmwmhxKLTai18lrNu6ofU
jSRF6k6AozUjT6CxukmOxny2CWX296HSU3zBsdz0vjgHKpdse/E4Gac5cFJb1tZP7syuDGaPcDsi
7uiJUhekA73V8VVt2ybCCtw5uHEMxZ/mcpmQBOCMLwcvFD51Fc5eAeYolRH6NvveVbrL3xA6+5ij
xog+jsp8ALtG7F7TCIGgXH23q4THCwmaTDeGDAlOq7TFUkA2/M6VzI3W186U0iW2jwiwLAOiukn7
Q+A8iFj3Gkii9wg1EUJK9rkq9xYeMGVBsRmh99HteBPVr46Bd2eNsyliK2tcjkXm8Yor3YfzJOpG
pv7Nhc07ht8izGLMCoeG9kxCj5yrDFFhhlcy4D6w13FQVTowwrORx5nIAadVDod9O3XEuvR7l4S0
VPD7UEJwyWEFIJIDSB1nE85dtJRjKwrEfhBBmlNgWmNUWeTwjXlUJOiiCIIZkc2/Z0gSMLys6BEI
JKm6uo4BzrnAmb+PUH8xbFoknTJ3Tk/tEFMDCRxSPXSCcf9ALQvLHgL/KKSkOWA1xvM7NHy/0xBh
mFjCo7+3E5M8eCwBnCH+nqXf2lw/flpaZfSnFT9/HXFZzi9NwWUhhYzQlXW9vUWNdREVS4V8+BgG
GzaFPBEY3QEKazBvxdO/ALsVMcjyy5cPTNac+AlNJOqESkN/qAQpQ7bP0rO9LE6G/V8UVxE3LvWO
r3h5ooRcR+UIsz2MnS4uIk/GBBkcHc+YK9u39yERzH5HBi8E7U9mi+bTbE/cWIP6CpvWDRNppkId
hIdRz7MM+RHF4XdoPz4uZIhxsV4lQb/fs9XeZ3KXRxigMPpJ2oxlGWin/Q0t6sHx42vcLwiz/UdK
15BALvw7ITMD2e/NLgj0+DqzpjaIB0rJde934zy8YXIyo4JODIJgs2X6WgGwAJ0VtOKh18vH/SGT
wglEDw5uIfX4ysJUsBNCeFLvqbsqnsoMoW2WEfaYGeuCfAIXTSWm8XgQ3+m6rkTWJ+0sfe0qIUp+
4SudQSLzFFoIO3qTXAmISB7kLqAncuQ4VbgyvmSBGyyJT664fo3gJIOivGaVuB7LlEJaOU91rY3V
TgP+3hgTbDgbTevi/AaansdVoMtOe4H6pmxnHPnBS4FzfDoaPfY/1AeEIots74AvFq0MjLF+YE+i
1ve4Vv83tihV3RVxn5SB2pBCl4yH45kwFOQlAsevanf6MtFH6epzCYr39i83U5kNyrKJ1sEhoind
47FK9uCGbh4NJKhuVLk56I32dn5liq+iF0nVWzr86gKD/nkUAbsj22+4CCWqHpx4tmI/7iHk3qI0
Ij/vG6gZNv+GfqnOHWU5Y7UkGCU1k8xsG3EETqKGIet+0Kc/86Z9lfmps/jVh6lrUsniUPQLpX9D
6ajM7QnuaYdVebaq2gWv7zUN43HfvshXdYKAjrcKcgKcX8be/dyvak4ThcQmvwenvrst/yhVck3x
BdfpkKE51/5jYlWv/hUPJXDSteieS4Ju7c8MJp18XiDOuPnjkb+gV0Q8WT2DXsTZrmkdcJ8ItlP+
bhY1A2XI2qxEouXvkvALAK+p9GQoo5U/H+IfYlqccu7TIndSOu8NIyoogGy6nVAXepwIL8Q6g7JD
i0Yc8VLUIVAsV/+8Ey1Vap3rbko78+bQygo8KCVPxqBYShXzPWierey9ZbOvhDEaiaW3xujZslOI
qGEb27nlDZnHmjzQ+pi8wZz01HguO0OqoxeTr8FL6Fp5bXULGv0tG9APD0Rb/OoHFUJgmC/aicHx
AtzhBHUHYPygtAADRIGQSQwXhSF9pAWIhNswqQIDmrXzVz2hzuG0mA+m7S3uSr5Mz1uJistQWy2k
m18mNJm9Aw4E6gUrzmU4G0j7j0kPxXtPlbI1RWZ0DNZrnuTd9nqLBNz2cUHYNmTDCbPuQOuOqWbM
c7pImp/Xgf8eQrmyt9m39mCSDSHp7CMsEnGT5KZ/KwjCidHegFNNmKQkAZhpMbhqp+bjrNRJveEd
FQxvWD3q3Jo3IkmTnVxVqG/Oci+XEQf6w7xD8HqkVWS30wATNDzA/1K4UJYWj50ipvBvyzYIZY+I
1nKZnrz45GqOvAtS+nqcJSuJ1Tfa7QptTjKkrN8PUwwhmjVSxuDtpH+YjedU9HjjRO/CA/AVUpfQ
HdgRelK1D5gbYQd7BT+1TOBaNDeBrAqmwVx6BCF4ycvro5HhtyAkgCOmiAyNQT69+wiAxxa8Payb
nOKuzw0txxzEua+rITkyzPqfvjDWXXTBGzuj+tAQO05t4XwNVP8pIlxm3x8VHsV/k1YlNO/99PXO
/SVBZOaRadJMG/ISwpduiFsSN+JUV9u/AvWOzt8QgG7nYs+O1PWdp5rHWJaK7qVVbPO4nH13KEUm
5wQR5Ol3D6YgB6pZGe8dCX6rVJnZH7dMWHPgIqROqkyx9lSjRa4ODYFhyOx0CgCaD5iz4wSjSnkC
p/eFNNZRTE2+KxZz0OOwhuoAJ+wydDx1hFoBSPNoVgK2gI8QdAV90Qnj/Np8tTkxPrHAe6BSDsv/
WnEr0yJTPq/xncBnmHxqFNPpR8Cce/YXeGdB7ZRFsDUJn4P6Yb+8gNW2DL8O4toDkzxnOGCwD6M9
sacD8lv/Xwmc7SPB/altIjXIPJj177dP6t1qjx7LFt0tKlFJ9eoSDetbx2sJuphajouFggLPmDmD
A7MqBSiCw7aXHDgw9o/42AD8rj5XNY9Kq6pLYKxPysHaESC130+7poDUKtr8kpGE+OjZqNTzOTB1
KUOJb4yh3hn50IJ6bdNkMtUUCS4NvxQcrVT/+KKiegZtmBYenScsYoH3CrR3xfuJgz0gqx3hXpeY
sKESHHPn1VrcTDkTUHMzBb+WRDfKmUbzE8Tg/t8qcuUAwCRP/y51CSrzc9mXtZgOgh5gxhXVgnAT
PHYRWRqR54txSuF/IcLbKn7wfGWFfJfavQTbbDQnAgtygNWPDEh4rbEF6M//yxMxCQPsaNOZYZHX
0/fJGcxYESSx308McILKCWmlrVCkJukfm9SXLN+lc1kaNYVL/q1TvH+Hd3AHYYEy5m1ym17VUs2+
9Fq/btuMflChRSJu6SAyzwavJRMvHNjgJhBxm6BNMEAFpTlKPb3ZLMUeFSIKD58yqL+96cDoJEq4
AIQN06S3Y9xiFeCFB/ijbSQ+FuhMYJI/9DySUEDW5Vm9sLoVHvB4JCGZK7jc0QfY5Gv4jvT2VSzQ
cyhMIUSGm2QnZF5Wb+UQPVd3LYcK0vvDqArZ03tSC6hKKCPSIuTo831XKjt4pPKn0nxoaYrymbZp
GyMmcbVL9SuD2UJcz8tsXYopnHWY0ZsoISJDFh4f117yJjc2EwcpuEEQ5LJJvSEf54Cl2dZeOpp1
QuWGir1yC6ajEunojmpbK2qELBopuc4K9XHfHq91FNmPSezTb4VMVRKorK8Yyqzl02Yjp3RVqwj8
a/v2zqUSLhyEIEYU8nfVr9ZLJ32DhiBwz75pWZEJAtv/CnZWh0LqAd7a3c9ixQB4jUOAarSjk+fg
nrCX5mXyGXdsWe0iEt/Jtqs61p9J/qp7eEW4WU+EbzoFFtnfXtRn3KkuiWqQuBs3PfQR7RnI67gQ
eVkc8kPRgIHXW+I13waixfZO7iIr3WBTgyGgqoO48+NVdwuWyhALL7+yurxOG5mzu79nC8kGcv4+
SNsl8Kh7fVkvcIzp6x2Q7hcLtoOjHDFFElReyLLxDhhmKrEUBAP3gZEfGhQ7kaoqzHN02VH7U5ja
haBnydPMxS5rjYb7p06KKmr74iRwHQnPSz/XlXXTL22WOOUozBrX0Mwfl3+mWd7ew3gdMrDO15ER
2Lgay15AnAvMo+N5u5Dm0ZqYtvHsSx+fPRtFQUgyJGxU2Vf5tB5fMEJfzhsdf6ojH0kaLTg8+wfP
OA3WpNiVtP7OpXKTYR1G/9cEaRpQcZDqpAlsI7tDVFwrOQrHzr60xMSYJqkUP1iLP0UOo7goVmRv
rGKZZNtqURXUNzmzKoLuSavSSGpIZNiSoB77VGtnYLNA3Kv+FVTrI5KO6DEKcjlxs7jLPFMELjvK
uh6Jjp/1oFzd8Aw1J19uknj6MecdhqJDY864wkH+KAd6ExQBA6+/goG4L0Y6jBJ7dlc7Dm5XILVz
4XVFdnuKSBbHN1yisSPXwv4WK/iOAHHA+whQJoRvbyGFclSLt+2QiL6EKJExO5pepZksTcFmZCT7
Wtfil5xjI5addvolZCMDbBap/tPrH7m/IXzmzKd+0skcY3qyqYrz+HV4mCA8xj2Uk83/aeL9ITtY
lww6S6zA8es2p3cNLeyVn3AzxFCp4m3DogJ/0qmBccUERI5uADIELL/WE/GDNhDQ5dbGLJrjp+MM
EL+hkwGjbNiP8XKcKK3NxI4YlHlYXJBAQusJFmnk0WmXlaaByVUPVUy+Vbee3cSIRumsfWHOWyRl
3ilwFOP71OPYQNKp4ik/Tm5kld4ZBAiDEBXU2HG7rtY961IL2VLhjCjMJYFfSDkGktaOOsMIamwa
PpTkdH5BOXkI5YsnyPBByzbk7gGY9KB38nAcTQdfNJreezmm6onmS90E5d+d5Qgo5Tb+f5HPewl8
PlvMFQEpF0tGdc/tzWpPS6uyOPh6Ju87046EpmK9ttQ4JCJHOHdX2F7Dn3z+Jj+INozp4l7jWYhf
NdiLudjepTIPRUO3L/j9RwTx6kDHzkEJLuD/64w0080jsywdHoPZ0NNy+vpAwPg958UFEfZP1e76
vODjNtvP+93np3DjSjsvxG9iQmQUTV/7SrCxMQhnLN0hNGoKBUi8aujKzaZStmW7xO2HFv4eu2jy
nd8JtaZdt2bKTB1PAPUF/hNLFsMEB7kToRclCyc5KF6se/+M4s7Q8doNKOd7X2Zm0lufxaHFamb5
QVbwo+GujbOhGOr3PdSA7P6kLaNpGdnAM+ClirwTrWj4wJstr2vyTmgb8UqEpnalG35qjmLbWEFr
bZvdnJ9dCPrCtAuBEjxRMWjIl1zOVVxROg+q1d9dBM7X57a4LOK9dGbi546gleBTkLYIXD6yHF+S
CHSjm30i6i/DNeKErJyjhzIokaxtP6TiRu6CpdVyzDfHfVO71BXz5tkC+iuDTX+ht1jYgw84eQx7
6xmIEBhop22Lqdvt1+c5b04N2g9ijwe3/BkzEsKwmSCJrfTDqJnL/i+JyDCS4eK7BDaL349LLhds
khNhoQjBx4JzepGMYRqqf3x/1NBmazGgNgxNyZDdkmmM4yCd+yfNPYrPtBfg57IJDq19ktg8pYVN
M/pKq7cQ+Y4WFhOMH2Zew5q76xGZ/rbgzgrcfKbpbKqRUnmx9NLPsoi+NUFsjhov/9iO2k6PdQev
09B7SrE0u6d2loTMwSN5fgGWf9T7dMXsCLfZmTAhJb1UmBZ1u8xHsNHliqQnZwkLNQ7jDtvH2owk
NXJmLwHL9BINrcYOSR0rMMhxx8m/iJhx88A94DhRaDcm+mDCJWbjB6l0YPB/IJIexLWNXKTjptb6
GDDXnAkGUU4gTIGkbi6mLRYFvIR8gYnFmwySviNYsoRbKC074LUUT3UVWoiOZM0i1zipqJ4GqTyZ
ttzLzbehJUUaJzfBPvEb28kYmHId49oh493SULfl9ZeqhvPzzZ1CmYzkO2uCD3asjbEm5a2fGK/U
/h/mXIfXH1mfk1psV7g4iEKUBuhlFjbb/jn68tznqXQlj+i96Gfp2fBl1rkUXJFh/hVqcLAd600t
cElx8x10G9y1ey5gaReJHV6l/w9WwxJ+D7mnmhDKfN4WRvysd95mXytMxmMn0do8Jglb96r6vrS3
62UMJNreFo5XLNlpmE138DTQ9/2WIQpIjrHDu2pkQSC5zcBqAgU6HwjtiVxTCZllJe0IukjH/80y
z01x408NpG9DqbimuU13CMz/1Knf2jVcY96e7hmwRzfMh3WWk+F9jfrSKNkuMg0mWWFFoMYpEZhb
ysDlZmWhYHYz/vN0X4aQm/33OTo7goI2mBQ50PHec8DB1kjAp2vnYzQE6AaWE8lTYX79NhRfs2tD
G357gkKy2Q039mH1pDBu9RskrxA4Xwr8i7LzDMnav9ke3sob19HvafNmnrA5ExcWHZIqL1PhCVEq
JwO1mAO6fbxdkxsxhpfqWKTKbndaWNeQZ+3uKcG//2b19YlgIt5xC5D5Yt69iwfubDD1PBQJgVPW
xV+Vki4YTa8VPCxAGAQUTCVUvp/rmh9chBNnNq4AMAWoy/eShTemxmYqedBmQKdPom0fZQJjtqTE
q2AYDjfjrMX/Ye5UG9PQIXM+a5ks2j+0TytxcEYKLy++m0O/yEJW8S3Z7yFrN4f6hdK3Ub7Duy6R
5Pz7o7FzkCTk/KHuN7ZZR9y4HhfAa1GUe/Q3MjI9FitXFxrbV4LQpqtQsZahpUaS0CNafalNU5r7
XF4t3MwlTaOT2qLwEI1vJoVl3ah988Ugajm9Y3GOy4eEn0PM9d/hvuJOdGpby4UpWnJaljcWIhRk
Kl5MqcVqYcS4hFiBiuF+vMwyTe1HGI3Zc1A5Xegj9oM/I97nWBkUTQwrBiX4kTIGdlu0JXxn+qQV
3JnkerBuM+vGxZBcPAuiptE3X6k0DiTnC3nhSCZnyFi1jbgfElotfM4/ISLVRt7trf+J0HoofeUk
VBB8QpqoxNLWpTeJcH/d6NVN1Vg81nn2Y+29GJ1SupOSIveaGGhdFI7w7Yx0mtBcBc4oF6Qgm0RR
far+3TtMBgabYmrhL1c9ouhLDvpOwIrtwQswRTj95JQL5s58lP8P8iJqxhduQ8vCMA0w0XIzhrwo
R/STRuHH2cnQGxZG+NcFhkmhwPCsggW7KQJoFqiosEolwZDol6s6va7GVGwOi0ghNBYGRAXOvlJU
yys3XGh6xtWqWkTAtfXfThFJ2LHS1jM6j2FDPh+jdIw31EXhAO+4I5zStTrLr/e+S4ngCei8+6Pw
LaSuWWuH6MOAGTSwCMbNlV/XHId5v1ST9wYil2B2e8UmMLB20mb7pM+fGxc51pD+wh4LGNZq5baA
ntUgY4RPoo3CJ5BV3Vhr25TNEIwrgJsGQvtTZ2hIw7tHO7Z10P87Cfm7QCzi3NsuK3Fh1AqHn+6T
tySdMsu4K3FpWx4Prja3af8LG8o6qHd2u9lcB5ir6Qa/+OZX5wYZaGPoqvDJ7j9quH2LE2/eNxwM
AK5vbugQUY3+pwlzkjsxRR4agU474gVclrwYnJria7tFZz+cvEPvHxwjBR6QgPQbf9NBGAh3RuXS
Ax5ICKf0K1sgXWmNpSPxOuHRTMPmQpwOKVyH34Cn8KLYxzD+OCbd/JdNIOuVxYMobk9xtQMKTAuG
R5O9vDwrRp8oyqprc4ESj4NzQIrqofDPkdeCdKGX2Sjy2PM76A1Mqoxakxwmbt2TOVNdnm/rzBK4
FNZQRwMRFuG7AQb13sic56XxJzhdmeMsDN0n5sJoU2vjPEDQkMTyPiXi3lSLkrCOyUH47vGaTezd
cW4z2hwPmkCvj4LEHYgz3XTPN1L4SIqi15/ZqFIgizNjUpNE/F/V+8vBCXc2A7IzwXz6/9xcvyTD
OPBC/9jkOTjW9SbPqK9JcUwEhNv6lV/dfHG3YXdDAYZQkEit+bUJ3JsJ85XOfenGOwRnKNFk1xD+
m+33xdhuR2ealYnXi6QI3E4/ZefLbnPuSl5bN5OQe4ofRVGF0/q1C77lXZwBR7RzpiAAT0pea63L
OMzGTlADUDaH7fjc+uv1zCuEe0KiXKO4mpADjnXYCUZ5Mshl1AFVYhzK59eJNowDTwRyEXnWsRz9
1d3rhVMpJt8saAeTZrHFTIdCzSZGOgp8rcPgob8Gc3P8OKktdt5jVbc4yTmQAaS72jyc49+FsiEH
9wiR3ePrm286jKvUnKjIbp0wS+GIbZzqXEpSH2KSnUQQK/B0KBCD+IEP1TnilmeyYOuzyLF7IkLD
Q0m6maCsI3+wchzAVq00fKvhPhxEJxmJ19W1bezHQXPqgQHcR981wb/b61HU12tKVxTamVQzljQ9
o7bc6QEZNLtsoq00YD8kamsOyKHEamP/yoAd8phEOIsInAeii58JTBtm23VQI7Y+uvCpNCVTlzQQ
dg6chjhujIloyk27co6A+m/UO3MIMs6WhOz7XJiypvQZiUd/T57WHE21Fo9Ml09dL45Eq7QoRj2k
l3AnayXjX90SrgWs3k5n3JRPzx33mgdwgo96/SNyPt1QGq9JEqN3DZ9m+4e+PL/YRZMglGne4l2X
sDuXoqkDt5otCo0xqcw5a5ULMYyMPm+0yvqXnTfth9AK0V6YNtyaz5sq8Gw0jxca09OWxUqJOUHC
yhjTU36gQSSUAiWIKP1OdkAxWF70QBohhbEIVb91SJEProGpIGFmFW1B+GZZ4hhejJVq4wGBgpS9
yeaiTCckDhtbxdgccN0+JiQaDvWq04n8hXk/mx/6f+H+LmM9iE42klvruvnbLqhWhMHpXQ3WtJv3
gDdCnTb3EjbHHTt4UH20IOIN1zWUElfVyI0oaeD7dZF+ZN76znsDhsVf0JlU5NJfYRPWXeS9K2vS
WMT/DThuFKNGtUTMD3DW1eofwhxmFto2sQX9eMDtNPX1L1gnE7/4s5jYW2ij87JhGIls4eltsDKd
xj/efVWNAcQcaqCfOe+XDOZZZ1uGfOx2DDmbazDtpZyPDm8WnJ7hdW+jBm3+NHMn0CqteDpl7Fi8
pYPn1YkFRj3to2Kz+wljghnM2wEl2XCPa43aJeQYmHmSt2DD8veEY6mdJpZKNVSYe4U/UvcxnOPO
OT/7kDsvzXwTRqFWMvCYT9xwcmbK5AS73jXNUIQ6ahXrljTJaPm+fU4Fy/6KNCpgKuLLkW/rwzhG
gRzOHASNCOOpBfu9e4By3760KZCUspBvoNnhqT3Ndh8qHP5onsSEO1Hb579YqLwgKzqOC9cji38L
pnjYHacGLCe/P3bloxApKlxDsLLjp7tfBUUHDjTICAGYOQ2mFxQfxAjDuAEJi3CdkMXsqtT0HUC8
y69U0VpkoYsFKcrC6oQyqQheitnuDUCDyv1JOlZ7czKOeB3RIpkFX+GV13T0L0PsYtIpFZBTONPL
+IgUOA2p33v+SMq/m02sCOm7HE9u1fwsO3cfIWwODXyxtvrBZh96gIhPiwtUXAsmLXccxXGF9aHR
i9eddMTUJO590CTWVvaF9Qp6cJN5SnLSScpQgASKIg8uQnubNZ0B7j6PsExJ6aR54vQzeoPv47yX
A0h3kv1JZlX8sMD9w6j3jx2f8j3eL11+VAeocFQoBH5YyOuCVoOKEr3AIlk+19uV62c3Pice65ng
OLP6TNpeEG7qDxwL1CxJT/YOCVvkDQIo5x/3rtQDZTtz5Ak9Zf2bYIcYaOVcyKDe+T+7VNkCoWsw
cY9rr+4DvDjJptLSXWdqZX1T2F5h8rSGg+GgNczumRtxiMSOryJy8byh9py1FmrQZTVun+R+stlK
2FW3BcrjGscuLxVaZalvSJjaK53jDF/A4fq+gcQ6Rcl1XtY1r2FnCxEfVJ88bbD0FZM3vkQgqDH3
oHysglqtO7CDPvaL5b17NGOK38KFyXYPQZSdPEmNNqPyhjIamp9buG3kIvufbldirM0e/9xqvvQX
2mTgtjckrwDa3zMms+Dj7CjfSDd+awjoW2DXfMIQQdEwDfK7pUdsf3UeHNUidEPAmEB2aVDVSaoS
vFalR5uEE9/Dl1IG7FyyPqO22EGvykXP7JcxAs4TCSp8w7fmjaupwnL+gvFnk2crx6zqMvjZKZeB
MVdt9mM/iQqtObgw0NBFQywl2NFEatJmc9XyF2tMK5nCJZTMYY1cx+MVplLBDdipDubFqsYYKNI+
ZJ2sIYxbKRWMYdG6y3lMLd9Gsh+ANjTJBMW/Gl22ImCW2mRNzyZKzWwVcTj1bvq4dMzYsv9EaMRi
Yayj+OWk/mCCKEKFWTZIcSBudk/V0p2xWeO8RIEmZMPmmw87uyudtW9QK0ncSG38PARq3YB7LVj+
Iu96aRecVDKvR2Bv8vXhrGFjivMomRyHRfCxqnpthmd75nwGGJoYnBsDhgcwWpZypHKpIeEibPoQ
H2oDarVgCkcg4dmg1m3WMInZiSJziGF3tNtuqtcDELPh+wD93M+GirQLqRFP7Uvv5AL6ku1GPK3Y
ic5OcPjA4chDbuMKACQq92USrS+gx4+G6cYTfP5UmF9WOwVUtTRBqs4d1M+YdxS9LY9jzAar5VD9
e5Nmr8uKT/Wh/fb4mYFMS0cHJ93NlQsgm+DoSuSjuvHZ8BIRoc/yJwGwV4uEtcqDz8smfaf3yOVz
eOXSyVu2zPTMKuqTcJeSEd9Qa1+fQY5OLGjgVzDyQzpP1jI56hA0t+i2XUOawUr3fhD4twn4W8XR
OM+3VzwRBQE34emsPUFdmUc5aLTQljUavlx22jhc29gnkk6CLH8pgi21cpa4hlRSM0Aem74tv3MS
UsKZ5nt+D20omrNENjgz9U/uawSw8c30S524ZXQpPMx2AVXqCKsOaTkszE6UQL5hHQtOl3LNGTxE
4WMsRea6YE5EFw5J51zSuv87Z7PHSM40OrVpwZPL2fm2rUVcNqDsOApuERFkCHGsShURhXFtHsvU
UGmC1huXKfSYDwvmPTDQka/9KSwNQgJwnOHhBEU6SrL7tkseFQxgMJbGueSKW2LUsTD4SxvZJ3Ny
+W6p3uTvnxycrSMSM15Ifma7CLB1zOFvBxkb+yoMgZJ1JxU5HCGn/pt9inbSv09spIDhJhE5e+fH
FEbXBac1v4LIzJO9uSXoNfWrqiiiGhHLPMbQmZossIVejbE5hh76qAj0Z99KgRxlvOZY18zj+REy
G+yf7wWwhqQowCrxR/ZNXobm+pX5Ns5a6qKV2LjRWRQzRy6PyeYsnqod4OHKtSstF0uwxCVuaIik
06dobjbDdvTFYrUab0k05OuOPvbsz7xEAs23XAJ9/3WOOdsuKryMMD/WAyJ0PAKy0ceqIv9JN2Ds
i3M56r3d2T08KXWG4AIIL1UJGSDKgBiSfAV8MyvKMuACHcn8/ZJiH9JUgIOiJGeAM1qyGp11gQrU
sJFkXKtFIbiDkUkngo2LI6KN9fvGXV3WJ1AnT4yURtQ6VdH7Q2mWpY+FHr1dsQfup5DCDA74mhhP
bfAsB2+UsTterzWuv5btF/gzLo3mR9pSi/A5tcMHszFgSuMs1MMKDj5zOZuDPpR1113x6e2e1RSP
rP/3QkPOc0eaKStD4rau93ij6JPcB2dP60k75+BIka/SNEY3TmgAh5p/m1OxAou31/2dWnb0sNT/
AXDkKIgJdY3X+QOENPRhR0vH+GerFk8lOlSvv+/nOYApbP+xSTUVRQF5yCFBmru8hAxvLpPVToJE
/pUCOPGojxhZ94bRXkmwHB+BaKNsg0vDVmVd07sZAqN7qCl5bPiuQkIZR48DUCm0vN/mgPVRWjKS
ZVBWSS3N+3OEoYN8BZR3k518fBfX7NmCeH7tluWbg3nzcsB77dRNYyOTYAWWsesBcXD/y+BTsXxL
hadUXF4BSI7WUeiwoA3mmDnuqCXfcDQ7AZRTVGr+kWAUGYKHa27DYYpIdsOd9SYVoDTJXaKFso5h
2GcbKB8Re2PjwgRD0yoHTXP/urjGHNflUdtic4XPM+d0MCJYSH79Mxd/9JYp0mVDtXwiiEkbpPg0
HzLeeYbx3qg/civ55z8Wea6lJb4psqQWnEK0BfA55SJGp6A8F2etKnUDSKzSdbtTrR6Z4mmc07zu
t/zi0cQjjv4nra/8gILNhxC+XiRb8mzemj1b19Antz5TzAsf110Ih92g9SASdCcYZMcC7rT9gQeZ
qrmkERnKtWOlXivoBmIEFsSV1fmk7YutSJBEFNRBW4JmowrPDNHf595S22SJbilPAsLfJ0RE6Jqg
2OpTY9Y0geX30UGHv5WpeDFksCcIi2KD5BePn8JHDiDIqXcG2Wpg0GFZg2DoWHdRmDkro2qwdi3w
hAFyOzX7iq8V0/13n20p/Sd3Njd1QDrBKtY2cxw6EoyGnUaRdCccSFtaGAHNA/Y7f5AMp6ynpCPw
mQZEIyIi2tLan8A8on27FKYjNyKyxHISIRsEgIIr4nxoNcRXZJKgKJ66fMvsStCLjUq1g1xqIDSg
Kyezo16jKzy6JoMd1Llq96Z68wjascBFK/79BgpRV+HmAasFKs/pzZIpMzc+g89SH8SHJ2QdunDm
wyKrm4e4eQuvVZh1nNYDt3XpG3V13cGd4Ffa4z14d8/43dYG16Aydwo70xKnZVlzMU5cb4KiJk8x
ly2wF8/DxlMo3V5qyiFI9DpOT0FL4MPjuqiOg8HT2RQNmeZO0KO35Kh0MsSUlmKYTo0Y0DhKOqlB
zAhfRPfRwWBVXITsbmsrNXSHkcj9dGPwGNfW+RqkxGRfNnc+NE2uUrFgskJP+vcw68483AZhCcGn
zC2NGgjwNlxgAFtbR+EWmizV/NfhQTZshL/7CKeNz4UC5+tR/zvp4ry0tLBXHG7/zfVlXO2Tp7db
AyULJRcKT3JnH1OT2lmrBduVKT8NazlqloJoslauf2K1HJpbS4yNkrjrtkYxH0xTF63N8OpPeSS2
dKA8IjbJiscqIo7+vKg2OonTj7MHprZto9JZSY0b3KNvc6Mj7dJ2FmuHY5N4FMYhi2ZXOK4UT0Y6
Lkho9eda4ea0v9f5s7JwZfMiYWtfhewcfHH/6mOIvZ3c1wFMYpdn3IkBpzMeGDKYAjYf/4KksotT
ieqvWjVzcEk22cXwkiG/SFK573eZeBwfzqPswRRSRf1mjfzbGZGcIqdmohA/Uw6r/LgSXGEV/Q2q
rWHJBaKVWLIbnHpH3SmD2Hco3jeKkrGsxqjg9KsfP7k29EP5xs8gLxvP2UAy7Htj76+YtcuIMrzw
mLpEBxKr/H2sFlncXJvGDCHisb+ISnWF0mDpIyGx0/968R411Sx8+iewGTcK6ElkGIPV7chpuS0X
D9X0cSyGq7++pwTveR5FIXlVZVg8+l58BRPDodxful1riMeSJeYcfgx8PJn6Od5kXyurm7kAvWGY
0gpM7y39cymsKRzQdNCGRAI1XrkOHOKXZZvjPI6uHDvhhhbtUFrWZimT5RCWDy4rX5S7kYJPMJIU
R3CMDGgfS3Q8/owIp6ttVmTXUqzyhmwjmLYgcUfIvMXyj2hyXPxPazxtl70aECPB8PbJf+wHZHbT
7o3HAq5U04NemeggpNdX/fA7UDrpXsDayC9Ut9o2aJ4VjeL6qExxbPYxoGACiUFoHMWB5WBnYssF
ICGYl5Gpn2DEB8NAMAyNnFtHiMXdy3AaRvffjLsyKqsQ8m9eAKKOO0kbH9tIiZ9awcuoPQQW7Wqn
tOFNjdQ9lUhNgbG7ZNbHxMuO0wmYDQdfXT7oAhAZwMBwx9wawKqt4u/39qbVaELQWv2nes0zFCKr
roAFk4OajJ0+gXgQVIAcAOd5T9f0F4hgDoIMSuLyvirRoHmDdEPkACB4A+vYEkH3pSVrQjK/hPMT
d99+dbWJemtAcZHoVaxI1DoykClmz98RdDF3McXe/a5sCqN+vbSjzZ83K++9rsJ6RarSOsr9oWWn
+vJD6GznVVLtw0L7lXmr0wI0slwPPkxxn3lw89EoibExCay9q1vcJQH3i2eWYLlYvGn/r1thphXO
ltQGjqMKwM+Xg0o4ZQDg3ZkA0IMHDwyooEoLNxW3GoM9xtlIRQG8OrU3n4n9JCEnkTCkS6izqonE
qRK5vNlCABwYuQJen3yuOIJT0ZO7+TWgeVEPhHosIfZgAr5VAk0NH+R9KIeAeSqeAVlh2+7RXUU9
R0jqTwVSqR/ZJFGTn8A/3dDWpOocuD1cT/cTaunNYFHN4il5tDSSd7S1b3PVbcy6iogAaDyUoSBo
0dviSjdPTqWYR34X3pDxGhSGw+6GrFvtXSquxi2ZgzDzAvs12BaUC5OnaU7nXq5gdhtfNGynEcY8
FcqpvckAOzjFVLpFAJdlX5f87PmB1EmMyF2uEr88oedd0RmDY+kp3s3wGh0eVl/heVoKIASRdL3f
EhlYUMZL/j3T2P4jB9QfQP64wgbeNuvmzWYXrN31OmmZgRZH/NxluICoZ3vp/new+a7D+EcFOw5X
j7TwSVBc1uzbtcW0OQdGXTXSZkvIZ0wvJiEWFzuAitxLWIVJmVVhSrYzg3ickAshhJihPJnR9Zlo
Xx4+v3uM2k5Tzkjv6O/8F1VUkJdFGUY/K5WDnGItW6ITC1QsA40GEjHVStN1Ca/zQkeMRvnomIGA
dmXsS4aD/H3+0DuJ+Ze+tkLbRY3OyJRUv6Jokm9c6GvjSZF1+4f7C7+TDRjzClygPj4cQs1LHKwo
wmZOUl+XKCOqm9TdKtcp0mrf8UoNHon5cyQHdQA0ypDX1Z3BwfJ/cRO3C++Irz2hkT9AHF/us20N
JcQTCPIkeB/EXeGMsbFjMjW0L83Z5fLFdpija5q7pTw7Z4D8xxxTXspnYaYQEgXJDEYp4r9drrGv
g0Ghu5hXfG18+XgKdHtfyHG1NULyXVHtBm/Aicfm8p9qqdbb6Vlqldb3KXPSS0HGuRCVl7ZOA/A/
TUwFIF26YOdUorMucnmQFCMyVlsxA0TxOFNJeafoSHeBbXKl3TdP3ezs06illNjGHC+WvodVV6Di
wvxDUvS/8R/JgB4MvkzwLRwa7nRjCHySmeexVl/zBuz+vnpUZcsiAcoOATl4eXsyu0IE36BxLNkJ
DX1vxnxYNqrHwfyvj++FmD4SV2ulgReltlFMNpD0yOZJaMMU07RhBFLsNVF9x5tOi79onfq1+Bbz
9ctrWouatVvmRH/BuPSwG6Aop5gkwvbhY4mGgA4eJQXhlOqLHc+4i9vrIMtByI0esZ6nLw7JNrXb
gNnKLAgXnYyb68wTcC0xZ1jT15joUzLPpsHR+jAbW1+PVp0oT4KAx/5L83KUrp4q6K7cRyQQmqXV
dFHqaGARbivCbX4bJbaD3+6hZJNxV24pUX2KvRu9MgWYW+SEofnAYXnuJw0Q3kA0bWPBdYksK5ma
z6cfoZDKqlJLkSFSzD8q9h/vvefoIUjnyRO6mRo9XvwPyoBy3CDZ/ie8TD17/ziRB5n3HKLC/h+Y
BGvs5dj3psYplxeUaIyMU1018wD3BVa9OfULHujAXT3Gtvtc0udhkuWXpsK/VTK6zFtNsSv2eTnx
AkP0fZoxHug/jHqdixmXi2w4OWZtXfUmnQbvIQPLSBccEGXzbVSgI0xsuyS9qORGuxHxxhGFTd5U
HtbiFtTAazN4k7dbeSHPi46Cxs/bpYYQW5mGL5AQSYtinzu/TQEF4WXbqoV7uiOZKFrlATbEdmA7
e0NdRqNZvuBptcHT6intao1+2Tbn/Y6PMyH7ghMUEmOo0OKNbycds14Vntf7emkC1Qv6BYfvTXlc
iPR8MF/dytIs3C6qzqIWZtY6mb6DhRZUYo889TLl8ZEWmPtU9FWr6+JOjzXhsc18zTRKXL/LtbeY
vBxi0jMyKtZlPG4lra1+61moEEnLc2N7RFDDV7VDV5Hy0QrLN2W9z1BbwJN3o8vjppDwBCa/mMEg
OfETW7/D8Vw1AGnJN+kL5K31LjP7S/WRBP8l6s+jelDyLrGAdal45Hhnz+aWaka+JD+8rGRvbeW5
0mitbALegcGuwEOKU2OXqwA+FLHTn/4FtDN6sAMOlmL5AN4NzVmRQld75HOWXen1LIPMIyHwpo7S
MM8N5maR5Ewnq52wftdPJ3AiL5R1oP0o4LIK40enyRhN/iW4JyYO3mtamvzCHzZrygcwoutumYEq
VqiQbT0iKdKggZ+tP4agTTqK59chfpE+Jf+uR7DwJ5xrxF0MATShqs2+128XHfXYrMXDAM4yPKgp
en+Ed37OKD0XG95UXKKp+Y4iPmsn5Rf+miUYqiop8g8E0GkobdET4RPoE280SDukO3dIKKweiGzS
jknbAalJFkuLv0wWjeOPmyLxlJhR0vjz7vItM/nHtKc7i004Ifg/Wo249iGB6irIPsLnfJxCz6xN
M/FJHgdOyKkhHuZzLD0UUKTEpuXjzEy/Hmer5KnSpMUusWhd6lgFrqw2dcNB5cXsDR6Mtd2FgqGD
o++Gt27Ik50kAj+EjhA9QMgOiQBUo6lENdxdX5on4JhOUbcZgywL9yPKiEa8hdHFrsjwp8qThJ0R
J1hn5snV9KxjyfVBJD1/H7ZK4mrnwGLh1fnss+ar5s91QHkHQ3oR5QLKb3673VWee8rkac3PNFZI
pH/AvbP8v8U1bdQ+PLJiwlmGw7H97AE9SLo6NKLqQ7pugEtSK8b6vgSR/NVqxXT3AzYW8GxYd/zX
m5QdPCoGQIActu4QyBiU21W6kdkoBcZVVXpwLdeQXR+fXmRZMnE96l9EdkpA+J0qd+aeoXh3yF6q
C1MU5b8mVKh86gM/Hrg2ofVaSWj6yoDF8lG0a4Gqk3kvshvLvvADGldeLS6iB6dEjAqex/txncc/
f3jWNz4R1crwNspPBAZ/mVOkjAaHXLAlgcCeLk60pdvhmwWOym2YfAi0Fn33HznyhGjQHwDZNWRM
OcMYfiUNAl+w8eGXSMszO/IJgksAr7UIELsPEEEETI0qFyKMw0Iln03ZwHfBu84FYGrHShucy6++
Rh8i3xCGjnQf/oPJ1A83uTS03EiQI/Z2GXaSACRsnxCAmN4dqmNnJVTxyDtPFgByNkrDiVvvtP5v
gbKFn0IMV+VGtYvnH1nJo4MpCPbsOvTu5/zcCrS673VSCr9VNH73TAp7Roy66yKOAUEYVm+Ba45M
oRiEfzP/vzlsfH/Z1E3G3zqnnkl56lsatsOTjLqhlEZ1turi5ipqgJceTw0YNIgJfYLEMqlRt4Th
ez1RWVwSjlueYTQNamLha8qeF84pCqBtm2UOYMpFgZdUw2ZYJdNnXIs2Vffqxigb2Wbcq9d8tdaf
3Bi7BIil3ZwN8dpkkcoQLdc1Uz9l+7f0Wwj6egHxevDJuJBuUxZNfs0gf966uvL5mKTy75B/dhco
QyJv2WWZkmNV+kK6gGffBbMymKF0IUenpzD67uQkwNNHH3IDlhwqQHvGP/VPNmeV81RbMeNDzscv
k4/jIlpkR5vRw3qSbm8gwKsX3wDb2XCg6mqH6XEejvx9Ptb4jURBbDIAlO53rF/isBSoNE/b8MGg
AD+HDlfKSkzsGMTT/rw6QIH2rHx3HOKFGuTjPN2v0BMV0cT8AUPEHZbxPnfsvD+C2qJMr3Sdeq1f
81ewnTW2M9U3k26byaCQaHlbZBNMqMdNsMoDDO9E/3xrGm1ZZK1hVt1Bv60QX9Ie+xnpeSJcHVrd
Ic6tZVhlCzDc6bWKe5XrRxOo+Ck9rIxzD6nDq0kCzKvSBpFpLKRBMebHwSvoIRNJliXJ6CIRiPZc
t89s033urnju/SDtctGHR5YpDo0q13+x7MbIZQQBVRNNqofwysvi/hCvd5rUSN+gsG6bPMxkUafl
6lSvAHt7/FfZEIbhulelLZuVJ/JToC6UVgaV/EP2UA4NM+uDqALmT5PkZQrphrQvUhUOYTmh/anD
8eQzx+P5u1UJgzXA/OpwZ9zhJEY/NIR5pd8TZnSuWveSCdBSsJXFdOQwbehhluczpKnDvHRaqTGk
ZIzooxUHi7zEBGLoan0AlewaTFYz9dn3mUcHg4Zno6HA8AzRqFRvsEMvyOU8eATQfIVJ/p+k8lFs
VIWE7ND0NwkTFsugNSVtkP7B0OlDhnYZFzcRAKA4TzTpSpTDw1w4uYuf4yBfRyINC2RdTmvFKidY
C5fD9vCB07THUf2tRz3ZnbPrIAyxMh9BbrIhw4aJAC7U0029LGEVhg8e7BVF2jNDukRBvNHlgcCR
W36lea573Glt+nnTId0Kh3R2YU9s+UWairqnFkyxF7wfqC/K+CPN+QAP/QURK+t6YGwvgkEq3n4K
/GUpbE2fVHTrnbkgdo5ITF9L50GjipEHHS1xWEvPGGoWPXBgP49ASFPVv1Dd7RgPcOd64hcyBuw0
5hrBW/ywrucmNBVyjrrL9LlEI/yGf37/7wuKb1cmXwTOIFlHWG3eyLUUXBsGKnI0jOLceWu3cgYq
KQK2SMsPicB18xN4WzQhmYeNbIJXodkN6egjeaPV6MmWn7ccFioHbEwR5GZo6LtpzlJUbUMeqX3+
HWvdpPQ1PTB9T3ZX9y7mIeOkgsauVd4TfKu/E40JTp0QcLnmcyVkBCuuziFyYtnZX9+cSuJwsxMj
zIxj6WeGoOEJ/UO3aFZqlzrQWrkRcBTl+vhptvxTOrMZAA626XkcXKpiKz7/wIEFUo/L8eexLTPK
7SKXtn+FdFfDVWQ9o/87GOKvA33rQZ2rjx3DRtkCEddaQ5Vh1g5g5kwP651kV4Q4Om7eFpVcQCUC
vTbj/spLvb3uDlox2u6pcDIPP4I+l9RZftYjjTyhmlrFBQvMau+5a/Gdi8LL0NI3Zy0Wrhdzh2/3
1XMo/uWZT+cYXiD3G2CHIhBSsmmeuxudq79BlR/ELlThVIitFpTpRw16XMarfGILIkpVWA+qeQpu
fk75E7hcCF2DX7BKx33QzLiX2QWUT7UU3SQ1mXX8BCveyJ9T/tmB7WeUHP7vxk7r5DCcgjbilduL
TMKxCfzIQzjtOPogBAryWFiQQRx7hDpfK27QSwiu2UxY2vO90HMtVMPAGbybXLNBUNw8ckVKDNG4
RcqD+3PdEGqChoJEl+HOZidDFW+45a7lcTMRNrhXXFb/a93l70T5UHAM3lDGPonVVLRwk1pTUPhA
9yQuzuH3ggHIxf2EPJxb7S4udlwK4gxV3U/bZzfTpe/bEn7YLKdNji/KeUEU2GoPvU30cgicZ1s3
Dr08HS7qd5yq/qMQrrWhohrcoFQcpeu48v9y4A9qmPT6fTBsJ7D6rYSwa57td2fuWnFveEtWX5hU
jLp4gWiP86hoGanRnzL205219wN2PqNZb/EQ+mw9FjpEoWGQd2/SaF+54Hyqlt01x0UfU/sFRGEu
X8nyFHWrj5/CZXMBDXUn5G3+B4fDbICpsb8I2f5h4HHeDlmd1E8eYLS6nFSOP2HrKsRPFetM4mHl
hON9HE6EO9cxSPPIe2/NSY81VDIF1tweOkYEe6QLmVvlu0ehEl6R5cN+XR/+lfIDG8cxldc7Bj7K
DOJr3AnlbTaA9YttCtp4nuzhnCD3oY59gMT8u3fEcQvMtiRv6uEI0xy0UOitCS6xLDCribpeZgL2
37BPnQ0aSTe7M6/r6d/+CCD3UJ/zDeQiFVzoXQcr79wJq1ec1irrfaNmS42cmnujAIkGkU9SVO79
b6gibEGdg72xDUo3bcuo3WZhn9Z0gh6Jbx1xR5rZDE2Sfx2lgJ5TNIK0fqFnlEqAmY3H182bttrt
lC+ZEldU/XmRrhiDGdvha33CbBL4MeACP+MXbNCo6499SwBA3ltKTRlyj6MEYb0kGjnpUDp4y2Vv
Y8+HNlfOoeNCvmmTidNJcJzTOFMHuEBlkopyNTwGW/rY3MFHwDgGbnv7PTwE5tnuN28dZ4HC40H9
oUnq6LtPDDwIOgOl0WjjzuCdl0JWwrfxYA2piPjiBaU6PLL1lVXRr1Ihaw07venBqozHuWjaaayA
4XDkFhzXXAJwK7E7RFxpgojmC2ZLQIiH3pVqjhjrfQiVMVnZtV59p9YYugifXv0tdhcw4BCazPuB
S6Cynlj+f+lWwQ7qpXYjaoZVIZPuVQRdVJ+Oq1JlpVRfrT9wk+k+wZwpA+x+srrTUjAfHXGQEGSf
yBHFeh/i5wsAI/eUjlb+kuHi0zP5rfogjD7rttqhu9N/DhfA+xrXCSuTVWCtDsFlPVHqpifVpHit
R3ME7goul+X4pzfyYfcdNMi6HtNLisG92ZyPvPmi67HIV2LNcIq+bmhpoZPRPLYYMu638+MWdkzN
p6w1/WmrkC8z8CX0co5WqWmQpLSaPYkYiE/KRP4Tcxw9FI4AXpvk+cgzOXVzm0nB8n1028UpScmm
JI5NIsdWHaYWd58iuIo3bx5W2uHoowc4pnqWbvpFCRMyuletGvSK1buENHPgaQD87tIeQCuYc+4a
EEXVvovKX8wVr81zA+da9wVaMW8lvNIhqM1wiZgvrOaVbvfqoVyTvp9++5Eic+pwT463fCV8+/tW
FMEx9tWzvj39UV4q1RyTbf6aLAaZNXlG6oFHmO1e55uPuBlpxEK+NrFQF3+P8wwEk7EYBEplVteS
Co4cehjEH+pE0TFN3i7bStKWCPtA0rZFA+sURUynK0yzIqXQshufKJLnJ3YzT9zoKjBx/nNqD2hw
Ma/66wN2cp/dJ2YP2rWeEhVUsAXrEX0alEwBUh4fMbLqb3CfiPW005tux+SyBmmf2NdY7FrkM3S9
3N+UH7W9+2JkFgGEBx8jiVlJfuI5hpNWtTj14CLh7QxKErBw1vFJ8xrJuO1yUiyRoWdHBWufgNQD
ylbECC4Vr6EfMK2vywY9hZeXrCYKynIZJNy304qi0tlA5MQEneNCsbUdflivtPxWwCCDgcSs7f/m
lT4lKMcOmd7kqC6q0u+7Di/ZTidlkSAmNMuqP7P/TDiiBu8x9gMWKJ27kMxwjs36k+N4fIGvzn/a
GnVQzU7E15wuQeNMZ5OrR84zEFDmyfUvhf+9Ufss3McciSN4jcskblZZuSRUkxJ6P3wVeUKe17t0
loZGDGFma4A//2lbvcl72JWrdCxXQTDpBm2TO+YBKMteWCK0nsQtHsVRH0v/nTLW61hsh9LDNvxz
AEqqsqll6qAzi0z6cf0h1L4lKxaAdm5oM7f98z5tMKI1mYT1QxE6AviFpwVY573Fj878zvQRSaZ4
BgfOVL3YqYEFSJ6oHfppu1K89CsNeib+kc5IdW6wDUneEqJHHMMc+EI8FT0JngAFThPQZSIRY1b3
JxLW/t5zjQxaF7WfKUwq7d4SKePtR6LSSv6jl8Ki1woPOkX2kRto1bBXIxUJIotrZEh5vgmQO6t4
64nxF88yHvg09BlxDlJIvQLBBjzXoV5k9zK+Uy7jApvc+CLAPrUp6IYqQ5UG4cbOeLXxlhUJz3wq
Lj/CXvOjCVA2kQFkuE7poYIDGrUsW+uNr20yPrTcwXWYXVrhsFGgedI+kG8D++4yD81NH/wVfCTt
bwnv6MqBXp+A45lWaOJnAnjL/SXzutuZ9QFtcwlKE/KZCl27uVxERpBGUBzzu2OO5+iJnU/iMPLH
FCpAPc7Buo+otG34hTeh9jKpjS10sH4vJvdMT2c2D1p2IytB+0qWodokFYq5LzPp2KLd0iSTEJ02
h0iJ1LNL2noxS+wTxxopOT9pukAjOF94rElR3O4iwdcxdtZmrZBV0T7ss1g+DLNcBTOLIMK9+IUq
OfzahQfb7vuEvYvNo+e4bB9xvI1vxmM9BdK3AgHripTTxzwU1gE3FxticE90PwXujGqQDYhuppvm
t2OKXW2mqwX2wWUUkSj+3XwrqwFdgb3JdodHiXJ/gu3tZ4PZUpD+2aMUgkDdUV2VL3M7TBFWG2x2
k1fV7O9+27lguXJe4riiBlNDRsBo8gYf/4kjVVoqR+GJ3U7kqyAJlOaTdrOTfXbMfdjEvjPTYq42
2/UUN2OeqdyvkkvZ+2N9GK4XPhYVCoBILh4EqOzgMbjv4OCVhH73hW+W8iF3KXAE389+fc9JkCkI
lxxWmYxXCl0mLu39Q65egk/PoOfX06P8975GiXxy51dEgQzm4cPdhS4N0zveEa2FNvn583DLe4dw
xP5l0v77eMmRJm2C3sVq5y0yaZmOCNL7sJgqa/tPUUlnBQw+Vu1A0rDA6RgWOLjzokzRwPqqgosW
I+I0ADGiq4FqIqmUgTZXkA2iV7nzMRgW/Qke6/z8W5pTUZvN1MjJYx86/Ms0se8HH6FqQqixUGQL
2lMuenTuVCMBRisSc143d157D/aWMnWJF6eujAr9ffjHhHnV6+LUFnPGgN9j1o9i17GXQDzJHWUQ
mPN7vYLxX6QDXq7YjQ1FhrcDt4mv5WIJ4U3bD2OR6vULZpA+RipKWz5AHaYSZXwCMMGSdG7TK2ao
JTB2IlyiSDRap3ncFJHSmQK5/228oGF+zq5W3g2EpWe6mnupqf2t5qhz6NOnewqdeaJi9wCrzvsF
xwS7y44HyfMNcG6jY4x9sGk5O/oNtuOxcfvjY9ilN3CclGu4RYpW7gIfrWvkRhLB6IPznXiFtQgn
YrDikCTAKXoDqGl7PABeqqJC22PIJkLag10f8aKxPPi/tQilUUetlqVRI4+PdFK75/1hcu/2ISB4
5OVbo95cBlV96J3h7B1uMMliX7Kmm1suKbzQj35fRDL3ZcSB1uSTQ7CbMn9gZlhGd2Y2d0fvXG6H
4FiSzCf7F0xEMPebVpyS44Zq0HSXLaOLAMDaEEaJ/HNIO9xdI3r/c+EcQ3d/Cs2lzOSQzBNM0nvb
wUX9SRbF/3n5ayqPKjDmw1iYFwmg6gvCSObziNXv3ScS6pL2U9Izqjaqeg9x9XInH5KqnwGtgrbl
j+Oa1oMpHEeLI6qvGp8WBoXZ0ErE4muMjGXD4JJr+Q3CrnXLfZ3c67sIo5VEvvQfbLo23dQfzHYU
9VdPdrjv3IWyxwXukW/+qKwFTk0HnyWiMlOhw1JtnitlBalg67v1yrxtBkewCLW21diEn13H2Y0j
/rH0i7LH7wTlGGlfZKg74omD2IdDzRztHLfViHbR/VgJQhHIVhs8lsvykZapFf7tPCDWz1H3vM3k
UgwVD8wnpEj10Q1TJdI9b9dlo5mlSwrX1EcxszJd44evpUPTgPIOj80gxYOq/qqIE1e2Gtfe92Q0
FuMV9JeI8gVoZQOxlC9a4hrSoSlQk9MVbufQiczFEYfed8zZr/lJdP0pTn+qPJ+PAqy66mGAz1KT
qQyzXHxbZsWlSm+iLvuOD2M+ZqFQkj4G+cca1oFWHAYkxrXUj8OYHL+9w++UqwVBmcsp/aRVtBtu
SJAHj7+VHl8idOeI0pJ87Ap16bH52N2TlxJncTkLnU4rjNXUbzlXbQ+fcGtU20fkeCHJAollAAyG
p894a0/QK8npWigbLnTrntvK77FKOeFeiwH7ephHNEXObBGrgCC40N+xD49lTuBfhH1+iRryFTXT
0cBeMXybWtfK8tn1CjUBBOoaMwh0yg41iWSc++BEAP5bLNLfaBtL8BQgz9HUmiAxvi7aH/lO+GiK
ScE/zOUYOPKzyPoj9c5V1BOMv/supPUZGHLVDIuepz3uvxJpfTlInBumSLJvLHbd6pcluWspbLGg
4qi4dp1ZhN6sNe27dWf7BjEcPFPioNRuMVqVEahH8wyGLF+vMm21rkMvYLG6BujDAJalZ0K6nOf1
q1lQyQ6ZsdUxMhA4ow/ZYAKJYnQD3wX694Mlb90jeMlX1bxLXN+gkWAPXuRh6zNCKe22HEIMBOi7
jYpPgnELB1SoQGjXfgiQGtjgctoqKoOWo+PSBJiI/ROLfpgACrvom3ZSZIgxcSpvf5YCSOySfLD6
nMEWWlEM5Dnj8ftMMt2fOcNKUZ7ykTxURWoD5joSnOfZx85owPKkrLdEC1QN+7oBvLvkqiEAHaS8
P8NE4e5GUM/6BHeGeyxaf8+YrIbb+xGMMDF2HLTixOi5JcbNLEaSehg8g171LJe+LLzMQMS9D9a8
WxvD4Blf1mg744iT3qsZR/51AHObVC9VPV6aaongqbZEEwBKT9dzoMaIrZa5BQNhIK5H0dtfQNnR
Gi0A8pkA7EM1WR9/QiO+N1CJIs8uHKE2uljFdbmSlcAAXh5OphKKzO7dI9fhU7Dpm9gdLX9ZSugd
HQbeeCDdaqp67vDghuJEiBGqRTriaaY1niv8HNmv5lz5TceXbOPH+ZSD+FCNzZcA2NPUy9au6K+v
6rHQVGcLN9bKLw/PxR/Pxj14T4X4gHN5hQqCJcc0Vm08aBmNzL29YmGBKZL7sN535ephmR6LaKPK
J8bSI4YopVdxSz8je1m900UleTysYmnAp3PqhVscIV4PK10WH7rvoZV/zYRKNaHSzyOX28h9gL1N
KfKnl/MjPAsL6ThS1XN63F51KqMKZ2juGMti+GuiaRV+Z3fJ6WOIOObJTpzfB9YsGyOH8KYMX/WF
mm6Rbb6YD+xo6F+sjpq26zAYawyDuKHNaAroWWDOAVMKkJmptJEZ4LjdSS+/ciPHBwSMCXVOkEWR
ZEV1qNNpSDc5Nh9LsrEmSeisXH5mxUKCgs3ltSTKJlOA+quARtnwhbfZVa/I2yfzlaMRhiLl05da
7rRZftz4O/rUJJKH/7wNneMdfwTKXgDEhUK9qkNABF0OST8n7p/NlS5/Xd4jqVtykb/dgtZ98jFi
bSdWXw8daUSYCHtG70HNLMxrLm0Ga2d6QXdBaISVWmLTPDlBrIZMsG2F8jfzgLw9yBFBQK4VuMSU
BJwlbhFETIFHTGC8v/5dVyDt6bTon38/Xmm2d9iVhMhRxvKue2hfm0jkmnA+eD/HKpwHbj0gB8p0
tEvAN/I+F9buQHetYYxmadamha4ARqSYe3SI5Q9t3WE3uq/yKR9edzbgmWHZC0JjuCWyWX0bBQhx
MLVZTjejVO7CbybCP2OPAgVr6WflZxm3W0t8rRXjLBOuDpILRkh2LbxqgeOljwZUdo//dXV16P/Z
mlSeaNAkdJFXcbVA82vJzg2wGcbx9GqQoutLBfcjCW8mvB6zJ95dd+aQIHQ8XWmJNCo8XhyL5h+J
rK2GK+vANfQVJ0Dte8U+u7QRTH8oxP5zrkclCTBmqWrAdlEjX8DFX7XtH26SCLO8YQBofQTpZ8Im
45nD4UzHah2nvgmg8Ke6Yr3IAZDJR+7o4bKyUsK1RtJpZpxOI/ZUVrHQYeBerUI+rXiF77bs+MHl
ie8AKgdRybPahyRv/39/tYJO9i3XikJyvzAAQauEpN3Kqjth9vKLriueO0wPj40KZT1vLCyGgzBK
Yx7GK06GCPIBWl4XUWlFnI4oYk2MABFsBUlO08jz42hJY02zZd2IfAsxzuOZn50SXHS9YkIGzbvi
jkXB8tSHWpkXg/T9YsYhbmPNIZ/cYPcOnO9qSF2R2cmY2yF1d5mIfsESQyeCytLXl/c6c3ZdkE91
OWcFy88MR1yKN+rg6ZN7Eg3/XvUSJd+RIlxdi5K1ztrScUFEqcvI1gA3By6IZAkuB0YWOEnGy6Pf
YYi4ixEE5YGT9FuXNxz5TCb/BlIclT2kFrQokzd4iQzAv1tA4WSK5ougkWyFj1EVd1RaWMm5NG39
X6JIqSxE6LHI8ZqOIclkqK1kBZIsJ65NnGFnjDcfgSTjYhlorBolTwYdQ7a5633bNUgdr2VTVERr
U+1fCWL4N2+AQBGSvBOA5LDt4KpBxVgft+GovxgRyr5jTl3tBBHz/Ah9ue7qk4rO0x4nGYp3zsYA
cvEJ4C4pzr6mL/Z4YTvP4G4b6Hk3lTy/fD80nuploP2xUW1ZSptzZQ2wjG7cZ7ZMWjU8tBF9sT2S
7LSxILrgqP3wQ/H5mEdRyIDM4rwks3xLHjfaXlmsSyuW7VgCjvwko24n4DcjYnZbuyogLeP9EDSN
QBfLxJFz4sunDThZHmfEmx/21zPNvoGyardFwYYCwgfu/l8HMTPZklFoijW/jX33opoAMPAsUefV
a2h6KLz9i07w0ecidjQzbyElTN8odf5WR0cD4WFvxxT/9qD1PBuR9FpelgFuVtxD/d3fUN6oMqyM
pPEUYpvMrwCFy3iosSP1v7H8g0K0jebbvNDNxcUWHawmKSMe1MqSxpP6jD/0O//Ycg4PS1N78usk
kC5HTB69pXYCNpyUbzrzu4zul+w5IqoS5VDuloN6I/2rtUzFtYF64HZbiw1IbWFZ5DqiMxdfkKzj
6XeQapTjuc262nJ2G7gl90Cxy6Za49ismfEdPq6PAJYCSbdHdCoGG4Q7r1FvYUIEp4B4bkuNDzw5
NMPszx7OjXiJufN7VaRB+yMaJKZBiYB55tg7YkQAvfyiWg32iWRzxqqxzukqppjd7LkdVF6AGuWM
GD9nmQIH33AcnLERjwvoMjUDMSKur+Dzend3U46IJaIToGVaCRcj7DqrbvRtUAxexO9qk/JIuRe1
W+ELRzfQ7THR7/JFdGAQTAak0hJXVhykJD00WT0tieD0Ph4CMclG07VvbT8ZLIMvmmOX1O4wXWnO
LuCWhmq+j0CRy4wPCVdVrw0qNWsAad7cW0SOZ+6XFFj8l/NttH6EMJE/OeGjkstBQMRkmfx/wF6t
+yyrRqZzXAvuYw3y5adyys60A/cCK1k7XKBU87Rn8oM1pI2szMBmS6TKln1xDePY0VtmOqntuH5E
MCtYqp0dTrDkCuPIFp6znHiwM7GgFBynL16Pp8GlJTETJ9lNtOVVCvvYkZTlkaoOF9IOZKonPsyN
N7FRybU/ObD5OmpgAi8bCDRUplWLa71Q7LkMV+l1zj8ewSuh+Sv2As2d5ntg0qjF7ub9Lyxn1HJg
M7OHROlNk3V+jYDKNwL9Zh3gCXh67ZxaOzq0S6zZdxsgJ+MPkiTj+NdIKEUZCuQ8gwayz5gBYUg4
l1PfIKyAiIWD9FkmFWwaTxzG237a/3Fc9aLwT+uLKotIynqwSnlco55JwcEQiKrI6dfkFXHdXk/H
GzsSazrwx+DnU0cdb4n8vGyMFS77JDP30VP145T/jdepxH+U03LgaldApIpnVrY0JtSziLUwwouD
lLgf55Dr5FXliDbdn3gc6bI442+c3wxRRZ3+WCi0lsIHZtpNlZh+KFn/+FweYhXrlN5ns6njNmq2
LTbhws9IcyxID5ZiV0L+hvJ++4xZsWRGevK258nbgwk7szftssWdFnpyGs62uh//oRognoRUkWLf
n1jpYLoMsVBs3YJZbC52dljhuG7sxnofbUJUlbRn/+wr3hJPVBanNl/JVKG9KwvX7pB6Sxrngsaw
7J2B9SAmH8dg73LOnJetTJ1kzNGMyvvc+T3tIOBRe6C7Vz2mfKsC3Z4bqGXJ5KEwi9KiA3yYbkES
HicEm3OejIXFVwB0HqfmIwsRF0gI8AaEoNaSQEnboen/neWTSWGlCBQQMd6qS4fMKL9vpqC/Nxlb
7jwgl1V+Tjj9T1oTMWeD/n0qetH5ml3hj2Uf/y94CJDISBSZ79Xz72rfapnc5g+kQ7GKc8bhkKpX
+0lURbFy8Z/gm34YebN+jHJ0eeg4jD6K18uw7a1faO7hRxaOEwd1Amp2TgZY4GdqOS/rfCQ4Z9eT
b71rwA6muvTZullS9b6c+BF2wq6oEE8Yt+HyEXYINTEUbMmz9QFSGd4uUOTSPiZ/EYsZyVwLwAds
jO4moEyxJKh8KJKJ3w+jHjiX5B4u5g8ZTuV7SfFg2EjA9+LTrTVd/Icaf7puIe3csgK/vIrIXmTG
1dY1HXPUZ1BcZhKQVcNBTecK0AolqLBotehk1zWM8thjXtT89Ls1gEGQI6JVf3TGR2GPk3+g428d
StwItPvEmJho/mTB1+peyNY0GAQBZrcqtjgdHSyatzVaaPIqPgIFKAwEOyuxdsUOQ8rOYJizF0CM
ZF5DBqg/yM8WHNTGur59no7inOYH9PLf4VNvSA7bCx2wt9nsd0AuLL38ze6sE0UruYDu0x6Hnolw
GELlxB0iPRpWSJ51lcJ716co8EwG8DbZLLFeVHfvUZHwFRJmmXtr+cfCUHE87Rwm3n/aRBKYDZAa
yw0JQAoWC9AVCPvGEkRtoeD0X5QwBY5YFYvoMI8wzzSnrEzkN4O7sZbmOD6GJ/CF2wR+MwqKvU/9
yHy0YQ4wrT1WRjyNYmLbPdJbMr0F7ePGfNp2YTzMbz/xTU3mj1TXFzLY+8flKwvGOi0V6HMN0zVe
G7xkm0hwZm69gVgzjWv3JhiQw37TGgwl3bC8I4ZTSn0uvwZL+sOLrS0FCIygtSfMMbTUvawTJKGd
HdR+fnf45owCTpZIhK8dcLXJQr4tDE0qp7c7erIrKSh1Wj6iGqahiKpJvWoaShsXK4qosxOmY+RM
skqnEgaCv1VA2qBrs5n4SBvDmUnce1Wa9kckeMdPvvhJ8ySKgEoWfszMpCr9CR/HGeR5QW+bVMhr
CpxOXZCAlRSiCEnkw21HA9BIlZAHez2Q/aYy5NjlNt5Vq6NTz5CgMj6UKY8E7dKCpj7Qk5Bl+1u3
74jIYPFVNZSrv8MkUvZWS8CcXfeMqGxjAJMdG3ZSNvBiLxuD5NXbmx5fh1RUlLG4pUSqWtgPFBs0
+8BcR7tSsexTVL3McOSZg7/8/2T84TNwjKpqJmT8Q9zkS8nIs9UCXnMB00W9Xvwww8AIBjXTYeFx
PweERRpoMZFpdiTcd6FLce2TRZfMtDrEgMfr8bBSZAYjZDqaOqLB2rRtcXz/IyFrTMRoREH3JTcs
IlZDc5TMPsB1Q+7Kx8pVFK+maS+Meqb1raa0CY/xOhIQyrjFKxqHMtl1tH1SkOXneF8tMuYfSEPM
0jKyx4EVo9EjYqUWsA1FyVvjoO6f9uRj79Y7Kv9pMjUiZ+plbHxUB3xpKvBUMZy1ASkZMXmkjwse
SrESlxJL8eTnJMs97dNbZgc0t5WKKK2oF1h/Ol3TrmtTnQxYql9Rh/kY8fziqcfSJnigPnZXiMSH
9wmarQczDeFI14c7I/SU6Tj7yMq5QvyCrOH91rYJAKKoMKbBXnnsnNXxbmp3l8/96l0MMrkWEU2l
4TxSj3ykKRxJQOAG1D5ZIH3a5VPe82EMsE/3phshDGS9vLXiPlaK3oZMUq81LDC/4S4Lf8BEPvEd
o2D8KACCLY1P6bW73IfPBwX/D4jpuX2bT1vzjJmq6THFF/1pQOD19FL5hWQ3xk73dEiOtg/KDVaN
3XuPNMGgfDz6/OWTxZBpgeAJlnKMCHYOIoCx6GKtP3YLcfo+Mj+x0GqZBeUBMo7VtOy4tjZeK5KX
6Q9V9e1Gs5OIiwvcdVkAXIE0RveLTFxLnY//V8/u14/unqd86b1+JctOIleJSXpAccWG/H4zEl2V
3JGmE/UxJRwztrkkvxVBlMT2yaNLj5PtNsY/04KLcvsmoPkU/qP0Sj8/sbPd1vMlKBx5ctpfvGLY
KIOAS1FEJhfqE1yt6XtxkAlsg7duQIzB0ADzFi9fCpokeDrwPuYFoqoD71RQdibdbjDh7L6VFDgg
eGWjpIxlSv9skbBBuv4KQYXLP5OkaeCnUSzyDlE46BevVT5a31ZieQFW7LQ5kemeIqmt0lHI0e2j
j11Uuh2IeiD5KJ0j0Bgn8Tp6Zdb4vq7M89FQsZvnA5YV0Jniw+0sOY2x3tA3Il19UJCvJnJr0ljO
zq55IM9OEToT+cXbxbARlAYpImw+FCvKNLxIH0wes++Hfh+b1h6L3Ovsg0/aVyaUwSBH3011Blw2
Tudny5vFHHXCwxrFNt6CpnGXMQFzgWo4XtpXJkd3/YKf3ccqD0S1gDp8cI2LFDHcJZ5x4i5aLCdo
PwQFvhd1lLjGTv0t/pW5aBQOk3D/TT0bnpMB8iONvB1AcmbxGRasA4lWQwVCpIbuwobfhyth2MoF
wW2DgswfqKD4eU5Df521s2XTofVtg81l2gtBwAagOISO4HXTqCSPE1K4oAjydImv/596ibXYg4c+
n09Crwq3PKEk/fuH41IoB57D3AOWNxHN227Kap0h1J9TnoZCyoAzoiNIQ/EqyZw2gu9wkGndfNYs
VHnZTGTtHHQc/yPAOjQk8PWFFufzl77UjVxVjCZucBTgRpINlyEjRp/LMHOSjPjK1Di9/pT5Vbvp
d9Gy+WpRD9CA0VRCT9K2Zh0OhH753WsTLGNvuhsUGpCKCx+T0Jcumaq77a9l/EiYNSDjFDKS76hn
Ix/bfbbq+h5XsGqGGsZ9OF1FDLpPpFQlPv3cHvNXsVNBeRf8I8IxrUn9ICCQZ/hblpr5sx/2JW3X
+PrWGCe0xLtMNUX7duw0rt0f6pA4Vexl3S36czMPZwc58QHVbCQqnLDYkvywGV10L6pYS5WR1sOt
Kel48Ni79a3oz5nPwwFyofBJdGZD43fA6IbVi/0cGhZTraIsc5KD0n1WPGpx1CzYt8TgY+4FjJPC
2cbyORR/DhBnusSekEk1XGr470qdwk6gaPSpdZ8A+xlaNlbX9Ofgncb2OjLk95QhI2VJk8ef2mHM
zxpLkEb+UN3oNpsS14nyeL4A0zvbx2QKAaG2cZ1IuQh3aHrsJ5bhnJ484wNCsII1F5x+M5kogv/X
9RG5L4xQyRC+gMGX4j6JGhcf+1qOcaXPJQ5BnBo4SkLpnCsqt3iUsO4Qp2ICUW91Y3sinxlAz2vB
jdU7y1miv/kNU99/Z3XywUuAOWZ9AnZer+BNOoFkTqWY3rpPu3xSj2PuHrzKjAu+hDWmEl3SEOHn
s1oV+yOhyBLZwFz0uNKHZNQRJRI0LiPAa+EfvmTbRJuHae32+DhRfJbHyMyG6CIddnlWoTsYAj5x
uTzg0V8OIN46OK2WDhb/wbpEwyetZS6EQRiSgfZlX6TjUATbElzFQaJf6cNaz3+9CN/6bmjTvmKU
+WV0qAbyvNdML1gOYovekIY2g5KjFso9f9CVT8wUF/Q60oe0QXlNylfGs+m/KOdkd8THeASqkEvF
V+61YWcmvPnWVuRGmZN8l1oHueY8nTDTk7sGLlS96viJcf0f8GQ5fY9u+3cGMHspLFSIB8/1nbIR
lyyTHpCtVNJw3fAJ5413J5KowjgGQu8PaPq6G6FhvVdGpePkJeIj8LdNbjojSnxsnwTNFN1ipMCu
TGI+eYxH6z89LaPpA0L/7/hA7eFJyLCQEZ145+B182zeMVfWV3s5Mr45CJQKZ/cokmpB7M90xsCC
aaY6arlTvdx0IOEXyO/fe/mh32nI4A4dHzRE895bbad+y1vGCXkvQjxtjaeW789mS/+f3TCkz5xK
LbjyLIbL3EbXRkGn3a0Z0E19dZfqvYBzxey5lDlG00hdWNd/PmGqQ8k9Z9UZB07LykebSNA90oR3
mEThBn7tEhZgiCFENDF931xHnZCis718nv1iKqh7FbJpkvQhdtW8xpYp0QrS9NRA0sO0eEZnLPxx
dfHj9bSXxLgcl1uVnNAkx/GGNXITFsBh2HiIFCKXLg6uGAvwSw1GK+V5qrZ9AAWE0B9sWlRXHxcJ
fh6njiBI6FJ9smO06tEz7DNXU86h0Y1oL50gqCZJAkN+AY3b+1PIdhCvsSP9ccb1bnTd8A60NWjy
Pi3RjTEVhFqNlVYaZDlwqDvcqfiLkciw2J8ewCAz/7xgLWI4rJBtcO2NiD291luUZvZ+/TyxJRL1
GNAHrT/XNXzQArK2/zsgCJG53WDaOQvOojhH+4t2lbQRsqG257atH6lL5dtio0drzEFaGkTnkDAJ
6qWjUjWHgHmTjsYxROUIuimtYQ2TwCQ6vJJgPXuH515zK0I9w38Rv3lxpAKsIfqkemLCd86AydQ5
g4g44jl0kXzEhOdmnpQ9J69M++HDp97btnyyYVbX8m4iOxkpLwx+YnCQl7p1NCggQgj3VhUqRK93
VS9kAjKJtIKw4bB5k5f/ZBKWoxIKtBGw+RdfsWzlhq7ZOQNTdfRWHgy6PMtz0VNmI7z70JRp0gEv
uKib6vny7URWtCmqR5qcW2ZR1cVpi55+DTmeI1wY9pH8zYRDHfCr7M1G/4BvprIDDBn15QxnP7+7
BXXa/M/El28snPBCTa0j5vMctzV5Bq90YgmFITTMr9ZMFv8t83slJtQsTlFJ2jhH5vqABp2AJ1oo
WrSxCZ8IBdJ4LI/qx3aXpe9Mj/m9Rb0gQHF3Ud/tZO8uqv/cWWLQm1BRolZudOJO5EHZ1WY2Km6u
gEuhFkKFcAJnmc/Em/qH/UYYrJMcd7ATf4FWJN6eY5o5KKYClTogZyZA8qem9uW0Mo1/I1cejgem
ZuAFh4/4r/YiL4cfpd28q48+tZXKcKTy+B1V8FCWfSYbaDf2yLNc5C3zthjViyUMjT1xbfG9KS8t
WWUjd1OfBoPJFsP6XkTLkInX1hACIAsOZk1natSiBuDXeCr2Hcrg9bv5n57nwplnh0JGwTvYxiWi
RD2Re1JErL4jZit3rSrZK6zWrg8hUaQ1ui7abBNixLw81wBN0u23TEVGoWMVeeJHUcuiq/Sa1zJL
zmlnPXliUfKXlq/rwYE4n++/8u+Z5rTUngmGcPCVCTqnIw0JeHie/i3Lse7ULWTloaEJ1TzbCEV3
8nuW0zU9kZ6p4IuyJbQM8HYf9ECfh8aVLOmwa2llRUvldqjBuTYHEi7l0ZwCEu/nFRdQGghfGKU8
lRqkUxsZ1hHcxYcrjNVib3jwatUR9/uTmOXX0ZpwG9x5ueIgM3pQi74+zzT7dQSl0j/d2K7wwWbz
LZ3onYXK9mGLj/Kt8B0/JDg0cDLuEX0dz9vOhQJOF80bIZgZ63CsT7ojBco5GY4lCWg34jNr/Z9N
cSHPbUKby2IzNbsqFglb+/YRclM59p4908zCX4hRbJdVkJvN3VlYuRSmzKK+0j5AwZUwct4b3nFs
COqb46OWJ2YbC9d9g466nZQ6zafjHb9NqpM6RpgQpEPZaqODVOXTVaS2Rl1fuGFh5uNZ+ZHqhAi9
V6A/xDBrYGrmgYikNo/U6x35fuNIvGkp/PC2/dOTILBH6OJ35g6nSraGPzRmPv8hrgX5m5vvl2h3
EfOK+rFfjIlBO2seVjH6a5dGU1v+faaBUxPTGmPPY90mkFnjFffpa19fq8ABIPAnIsSTn4ep7KAu
KkIC8I62W9EL/m5JhydQg+Y+uXpzP/DkyhsuAXPpmJH0vB1EUff6MQnxBQtGIfmBqYV2MNSMB/8z
mZhYOTJy7dM2qlcmmIVDNP1OKmco00f26YlmJaVsWAenm0Cd86r6g/r697IDpkgt/VZKW+8bRb2O
tjANQd1CvfrREoQdEp/fUEbDsbmHF8DJGHfMYvYXOmb9VRt65Z3YRKm3qQs9dWmLefMexNpHP1xR
Vhqsqn1K098nV8XwKKh+exzaj1l0Ifk2H1DzXyhnrDZjy+4aCYaTVxy3ZTzmmPLBcYyXSdgSJN9j
rdkEFKfnJk2X4kuJ8zhFqd5Sy0SUM8bWzGDcrvdba/Zi3I5GjCgYeMWtuFmqWgF15tU6MeVAMuzf
ykWSHJjDwD4VIFjjlEzsXkv+ZCBB5pfBHRxkJqJNbAKme3oWZGBFUfDW9huIFoCRAm9xveHTdxFZ
oPHLVprWfM1rxxlHkQ4zgR1J3lMm3CvGJrdk9qVmTa9iXKatuUgKwKt08T9KowAJZqyhccpUnTNV
oArJWJsTaUoHlPTW0NtX3Son9KIlgn1d6iyLqIiN1vBjnpA4WUOckAHubvYvQWfzuPmgms1GyqoO
w/r0klwdM3POsSymXVN43t7yJv3jfG5oinnCKj0fH0BCyn0VGQuH5U5vdkswN4Kw+seD5SzWoA+5
0Fjx2kyF4t44caCtmCQn51IB3bh9NTc5L8V2C/UVg+BZuSmS4acM7Pgmy95yBsapiceb4oZbpT19
ZCdmn+fwhkD7wSOaeOltFXxNaTty4HfIT4KPpVb7L1CBM0WUeqSSOtl1Kt81Q88xbkSkfaJrRZWh
6z+oJXGSGedGa5r5aC58pgn0yEB4v7DRX/DrAUTQp+Y23Ccz+c32F286PSvPOX4fAnIq2XmiQ7+K
8HuwG0fsDvzWwXnB6eyC+cgId+sGsf29TjjhKu0/1NDkbLi299GWy+HaYNZRGxib3gqUMOE1mVSy
Ikm3I44mMvjH5NWoHw9cJuNDVTRLrO2t8r5sqCm5ytTxN1LVq5mbdXoKHNGjPYE67x6qJqJg1Wyw
HkzKFuD5Udqy7JiXw41XPwJVhVKwIwydvsVtQm/JpwJ/K0IAo7afuhHIMTbEAwqmt+pFTJx2FyR2
EDj1D9vlOOlgNugFXa6y4tR9seQSU/pU3W33mDeB51fp0Mm5WRZpGensqSoeUw0z6CZ1gLyiVle5
C8+Ie0E0hVelsdnVJSOP1Y0SDWBJHNafIZsDpt521DwmpR9idKTfbkDbxol6H/0wW7zsLN/xYcSn
pCey1G9eQgzeKeatXr1syFO3g/GqaJOfZfR6krp/dMA1KwGmxX+87bQR8FVzR7R0uFlNSi+A7SMG
evVUIEylAgE3W0M1qX1LUxm5hiPwjLxnLk1Y1etK3UdI6BDLf9aH8Qud+9i/u14W2DszcsEgzVKk
j3C+0HYwNquQmLjBxPESXdMejsq1UZfKs6uasw1pNlWKw71KUVcK64IzPp1jUC84FHd1NCZeS6VW
KmR+a5T2fOYAOt4IJZOH5TcFOEcLhD0XAm3aeDnesjsKI40Y1Hz6EGOfupeyk9fStDVja/zVTuxz
hFFOkOJ4pGv+tGwRHdpJziGp+q4I879WXidFVVH61DZaRLII3UB8gJDfIrbyotxOUBE9NLiX6/IS
JZWDIFrwhGXfHySdT3A+K6YiWtYEY2Ktn7+X6l6PLJ2FRVAUBJ8wrSSZCb66tvOdwvhR8tFqpJKR
5djfWPkWoEHlxfiXxDY6cVw9rYmkJbSmxDw65VvGJV6xNb+4bs3vxhC7D/iMSindWeLaL8HsxBIR
kWTe+yaUBvAufQvaqtYPMxSvqELU6+HqvUF+Ik2beRUTNJFMOQ7sjschAI8mGEbQn5sbMNkY4LpP
Fks7gOc4iAWbx0pqGLx5cYJMELI2e2v4JasVC69Kg2EAtoUv15O9z6GDEf/wYex+atrtqdxscUZ+
Ny3a+9GnHOBrCHBxUEJeCnYp9wpo2CHBY9snZlnW4VPrPfwrYIU2i0EifuBuN9EzJVaqnhixPgSS
UkCzZZ1EtEtGpskOUyXY51Ww6NoRo1MCwpVGD/gF1Pu4aD1J7vhrtndhErq9L3AcKmWRD8GHctf5
fn5Mi6bwTxULTAzbNBCk2lWN85dQLNgvCFGXVZ/8TRH8BSBwQpRH5Evf3DyrLrGEI947lXRIc3fh
fIeLuSOXCA/WwzMhpSCuWOqrDhq60Eya92FxM5Xuh8hR6hm7VNc+6l526QBpDQt+gg+/bKDzfg8F
4OplEG/btjao1qYqUWqh6pvudSiw4JZANjNLcbFMwwn0ETrRwEfB6UKTGcx797FO5KxjcgTc5SJ9
Uug5uXdZZHjdW5/vdOFqHtoRbym3EAtPjLFoP20roDK0QmGiheNhPf5DNbu1IbOdhRDDYV/FgwvM
KgcRuqV5dRARj129NbrR0O9dRwgXrwunrwsccAsnjG63T0/4MAxgnW9vBa+TGln9IqjyiQ0xGeIs
k6cMNbkGdKWbMcxYlOrw7Vwa9HqS4/L97wfQEVd/xBE27VwdmaOjSpBuL41eAm7+nQ6f+q8P3WO4
KzY43z6QPH0w2Mnh1CwBJkhplgK+eQ8dIAwKvibCcOeMTmYejwlTHzOp7SoU+xXgxPPqlYlu63gE
ImwTLLakTPBmU0Yya/3HLbyjdYDLK1aha/Zwp183vmhvLRQ1nKAYQo/AE7vdscFIvfCbfYWt/Ex8
10LVCmEryxg/4DLw97pmQzzsp5Kvv4/wBXuHsTzuExX3OFWnhpv7HM6LwZ8v62DeopDUXQ7zpmWz
iQzcB/nDK0tcIiu9zz6uCPjK63v3cw4qPHMNStSeTrFtR7rHbj+teifSMBPNCMj+k6FEhsYBQary
nWqAPxs57gf0VcET734JagX9TeyiQ5JAUfjHgbNa6Qq7NMYfqY56C5VGBXhEBD76dzr0UW66dqG+
nVHgqI2dFyIMk9MPZWCQ7BZRE/Y3NGaBn5AuwWXwBzAUlIADEEbWKVEiKFqr1DbO/8lHJ9vMGg1/
cq3Iyeo7SP8YSzJdr57w18AZDIIL+vcM9SH49yUvOGZSWmcBplNfUjnpI+Mw5GI6rKdFekL4tmgh
sHJ4JdhiVJ4qOQTnUOJKWAW9N+QAzHarZbPD2Od96YL0vxoiVoVeCtp+FQST9n/SFU7cijZHFICm
wL1+rAecCkhKVsEMKW7bbn/eYQtaK1CRnmLk8PMSC8+gMLbQXHtSr43nDMI4qTtJrGknD481nAs5
Nl1itQenD4KUMeDtc76M9W58B4PudfUedhFjQcSGjPCq/jAtZwjo4eMgO74gYL/qqxEmvBso4/NZ
b+/zpdkyrwk+fs1NW7kqHoy1BIAnvu20Fg9veqkZ1odpelLMzpxsbmn3Xau/bPCHeLpKdVDqlaOE
UqfF907/xzHNuHL1o4jLCv4GR3pG6ntJ4mQtLH3WaHKBqwu7BXdMQrFIO8J/rNK5E+7VEX5+1Gjf
rlh5DZXqhDaoIHHotPPFUBd8tvQ8l0EsOXf+Z4KsT5nqGRKWtnCUlZuyi2Ooz8JtkK5sAYAf62p8
MTffhTXklp6frmMABrQe8NXSRVSjsam/UNkChWu2R2Fcsxr407PUtJOOKlL5+ryIISZP6xqOFiAd
O0Jy636NaRMv8oe/6m8GMvRt7Dq5zvMjwlAn/qHafTZq8unlYWXHDlVRQJISS70zK/XjriuprfsX
KfnNR/LLmec1sXjqDwIniqQSF2vt7Yjq7Zb1aPaaoErME41Zt6PiBbdqAVC6IwAxW2kai5MtA8rb
ok58/DJKUaOebPZo+uKrJOYoU+6bz1BUJyf0tN95bVoIjPnqa+2HtPMILvG8ZqAK0ch1sO8hj5am
XunptoxU8h3B4a9Oq2evM0fhK3JouSSJC+X5tbtGTrw2GH0xYt29dxnVKETf9WDXUn1cRpqwO8yQ
nErs13RbE+ItOMQJUbMxvnLGl8TC0Ov3iCbyfcxlJF7yvhcS0RwxR/hYxRg8b1xm6J18r3Q9p61F
oc5AyeuW1BtgP/qqIVnLtNLfJmZdc/8yqdTHj3Y8WDsSFnbAY1Gr2mQRr453Bp8VPfpasbFqsiyS
Mf7ur0/iHrV3k2QE5EtPTmTfi1dgciDh+TZ60xx7Jc9tN4eBgr/01esbSft4EIxuSJvehl3HowSI
65MsN0kmSLZPKIra60YlHe0iK+L3owaL/CgjN22lqr55f8WgLdbBUMvzDCmTepe7FqAfG9jDwS+Y
DJSQftpRPy239tugeia75SBmOEl5+KoM2kXp3zFq8E8anpNwMVtVpdi0LcfhElVUCnDbLSG+UIMB
wIaoFRI51PP3KrThwGsngmcm/htPP8q1ZNWT8k17dwuiBuP4m62y0M6qbDTKbHkHv5oUJKkMxqkV
UNjNdT0Rg5UYCQDrSbExU8Z9y4KlXA+tM5MC2uYfuWZ0Ws/aIJDOeAFN6uqJMbDX8/lfC1Uj7Y6k
F4Rw6mp3z7UcZ2Rk+CoxvLNssRkgMKtCT0UxJ31DYRjMzexrIzQDnLO3GtJf1z1x9BfLyx5jHOuA
+lRSbQsAzWkErP4tCyPJ6cxEcWZNIt405XIKY2h91GBYBRVTSazdRv90iPrvRDkFVB8PyuXsIKRK
ouI++qM7V4QLmZ9k07Ep3MUwMVf4H+XkrbPV/1faTgroieQzIjQI+j3wHQWvfmR++Ke0mBMPe0KF
zVkI4xLvU+Dt8FIRe1IgG00oAqeBAAJvxj3Sv0Z2LCjTkOToyX5RWMMNgVdNk37vMuZglI6eLe5M
N9ibrmQspRCD96eol721ULV82cYEq/BqKkTXUQG2FLU59RVrzqhrX1Q0PHOs9/yO0t7JSOwd77oz
JKlQmsAed+sIHryINgDYt3cSX0F3fsBIJLuB71K22KTEOEuY1p0cz0yEu4gUxsMxu4U7+LvJ8Y6H
RWVQ9zKettrn8ajq5ZL4ZsSQZzpr0bLoRPj4uLaGUWo4Lrw8R9sE0B2pP5Y20jdvlQBrST85o5ie
xmvkpCNeNrPSlBoRdnCfwrNzyvmPsKbHRntGxqWMXB0aYWXBxXbjKflarLYmPL32TH4CLpRdKyXS
TR/mxRwP+tzuy9Ps5Cch1BtbB/O/gaHwMSAl93bXDq9ftrbr+Hyb977XiP8aVMNokHn11lJ3fqAj
9FzrYp6JaJj/uDcW99gLwZeeKhR+E/mlBlxNVTSAb1vmwESO04pvbVSW/wuBbXnFvTrZKnxn8pNe
RbtK0l7+FOhU1f8TcGbHgMp08TGzthTIRpTrebE8YEwNrv+M7R+EaifIH6O/qhNn7kEVLBnu+ByS
LDbhu8fZbtK7HvBl6DS7GosOD9QNWEv7RkbG2Zoa2dP7Of/j+dkAfXH1jp+8tNdV63pOfSvvOQI0
3/tXiUEi8801VG46QEKywjgHHYvwEYDUIWIXfLDndOpyh69MRbd665QSJ0G5lUtk/KyBKltEvzlB
BAcxYzsmGx66VyvKCMuGgFl+/mKfOOKxHSrcO/7BvesyotIqS3CDy3WZZBMJN1d9aD/dirEOrVuV
gNls7NVyg56jAEHzOfj+zK0ppMWijb9gm3NReY5A7KbjtlTFy+AlTq2mQGfIul88yyGm/R2lplGG
JKkPhypGO0WrLV4dZZcaD2+pf+z+eN7Cw7qJ7Tf0CCKQh92+4Xrd0+kkcykcYLoYWJQIhqJf/MQT
pbb0T9AUVzNTU3lqWSjGtXbOROpurWdiz2gYaI91vTSW+etYf4TOH0s9hsyMRbnBeB/qHvJx9HE6
xi3WSA3xE6wGBXsHOcC18AldWwCu38U/tN1LRLeX7MsGMoXS/+GOfg7N/uzb91Fr+tLiR8Qpovl0
5lYSM9t8GA+kekLx+o5XPK5bAEJ197t0+7MRI8NXWVCx+dgkWUhRv5cnqwVe6ALt7fvdRk/a5a2H
T2u6HtGaoACiURtHKcxKKAQcLr7bzvsjHk3VSbBoq7alk7el8W1BcPajh+jjWAcm4astygMa4XkM
4y9Oro+qgO6vkyExbZrtoUfTD0THoaz882DPPqw9jTKVgJowAQ2vD8/jFs6KmOBmmBVV15VySChI
OllTxUzq9n+RYbvgubEQeur45n4sogjxls2DEu0KlXidB7vCgsdmYatRxIwrjwZGoD7kEaMUcroE
huuAK43S91+83dflOjTwMs7SeGCuN6IzOgiXqs66M3Ju8lTBO2DWFS7tAecfsjtlDsWG5vxvO2St
WlPM9WPYd6xwkMSicdInGIJ7Btp444EoKOTR8uOMxk6v2rPyTZTc77RuPHJ9hnaXI1i1TVjRsrTN
cCOxTqnAOOXmSnZGXDAJZxRM9qEqc8n3UHmgM+sWiGsJaUOMVeBWYOaidAZOt7B3nWTyRwpcX22x
wVQGoys7hPtx+2cCReW8iF2bnGEVEjXcU8/wARi4ZUAYPwARRX6PFJqe+t8pJ2rZslw3O2UsKVqt
4VKXijhjmVeDF2baX82AWrmyy65SEMdutIZGsQMTOwfPOyDoSQAGtmWL1Z2WHyzSKdvkR8g5iCf2
TQckC7jxVkD26AQJNt97Dl0OBqoTq0VWOoJFn5ZnV7kB/HvnjfIt6jQedzIajtD42PyXIqBl3h8u
0hvRgMgjBMu41XyKPvx30jlKVh/G8n444j278RUvTLIIghQ5FyPX5lopr/y/IdJsw195nvAl1I3F
akzXPg4AfMQB2Zpg3lcX5eNRMGIk3LGW/HLVm0Zk40aY6jeKXXWAudDFT/K8+b3Ug8fFcRQKtq+5
c4wsfR/1PO4POZ2FTgowRsmCDD9LEbYfP3nPjNGjGe6h2a5P2DFTWgMyFEP/dp8VVxxp8l4xXnHO
YFLr5iXlETPMEtwhhwfNS9yeCzm1JcPPzYCqXeNLkWtHAoxt96UOWOFZt7FIRvXv3dUcOzfEhY20
j4I8APfbSOozfKhcKaGyUVAgOHm+7ZIxj8RFW9x8kZh0IR2mgiOe+S5xHMyDypbMrzsNO26VXycO
Ix06tX8mOdCdeajlUUzbP07EIcBm+XpTMafFp5vNxCj5vopvplEIimxHFEDrGK12nWverSROqQ77
a+v2jS8YR2ivpmkA8NBepxz85mdQ7TUG9LMXiuJc4ssLmVahaMiNVXMWyr5sQgQ4K0c98qNTy7OZ
OlTtzYOZU9CfYBCbSqPH/kJfCq0O+NBWdXwre+BV/b+bLXmbYvl6t+ulYkKXGBqD02i18RFOGoci
972X3ukxZwGJ7ZwsL0cC0c0vFbLskzk7VlT0F1Z7MAT97tTgJuxlQlkoCuNRsOi+kuIKGZOuTgvX
86LbnMhnuvwfYBzQ3ulcK5XTzrHGWmNY+XXdGhwJ/yV5BwAL92SE0/NSvndff1hLLCZBcVw+7Uzp
1nOyjw/Na/Mgraldo74KuI17Jbq+03CIvtj42WYCDhrIaarNTmiGGolDDTgRu7HoxMTOrkXd0G77
azylmu7IkmUDZ/C8vhUHZW0LcKNYtG/CMPSe9L32kYE/JOJ3bP4RnkZS2Nhiizp4iXE9U0rr4ECu
9ElhfXOwK/4CABLV0PASD8kY2oYGfDF1gRuI6Poc6c0kXuSKPocyZW/xCkhckJJkRdU5UVspO30L
PAPGIPqtkICrynX2tW6ciM3/feG5mjZEC8LQ1bC+xD8mpp0J6iIWVwxSGUJG1TuisOldiIsOMUtl
lIHHVAf7cCRAqQNIo+dViwWdZ67pGWwj6wMqg2ZlDU4N2TYi720AIK96B6DXi9tlSuUKNDf/DyaS
otXLfY9vSaDO+kYidu1ZE5oTpEbX2a94I0mlV3xSNviHnyXJCQbFEIvQHDAzvTB6IzKlgdatZvxw
XCfxJc3hYMD7B+SXNLxH7vjW/dnqO+dRmYjZ0J5j7Q4Du64Gcqxs2VwmaXNmlvpJ6qItoZXnChpd
Jlg98Df0eR1QQD5MJ6usdEH6R5eKcV1uTlWx5InHLWAN0t3UnaEH9gsdUPT5THORAgvoemcHGH/t
oZuPbOBi7a/XCTpeh05IiEzK3ORriYNd85brhS7xqMyKm+z5KPsjZxmlfupteoxnm5q4h4NJBeJc
iD6eQw7P6ZUdSOght8fVw3rpgBXgh2ToXfSr2mLeUxck/wkpDNMXrol0obE2xBaVpMwGxj0tRtLE
zN/tH8rPPaHOM8zlqLsYao4fZpAPX9dQRnxJlizdWZXhpuOOBe+02fkg0jY0zeCsmTbrbE80ODR6
6EMIdVNNb+6LgNJbJGK8SzwRRItggZo3VsA+CPaSVxpPVn3Cu1/5yo0Zo1RDWZkEqI2YTgaHKsvb
LGVD0uolXvDgEsu4N6dVhNwsdQ6PQc+k4SxFxsp7n6OBkthmFmU9gNGeuYndSrEETIo1UeLMf7Ha
6D9rDgM12oMBILhDKaccukOpHb+rtxKqFHh5xdxIcUDblJhRug1Q9XtaD6NBnBV4sBcLHbuXHg+A
3kT3QocJ+hNl6ynPs2usPx8/Pa3rUh38yxTjvp+TSof/G3OlX0MVmUk7oKTwwNjE4z/8fcQRdVLQ
Pb8nb1Mx7ktpdX8YvgLM5nDjAPcUeif9b/+KMog4M39HynWADdGIcE/qu3B5uJv5ECqkjnLKUJNu
PAHHnIwUotnjpGffomGxECM/2MTTfGrg1gYfqPLZBrXOvRQFZwfW37OxrWRCZdiAIxKWp0h77gPZ
w2ggrfEC0ReUA5TCCM6zT6O96EEaAgm71ow2VBKVVATjiBHtrKo0RTZN5Z31uKX5cL7he4y0guFn
bKDQsu0Bvqzf8T6NOVeqW0fcgFn7aBQjw6X3BBZtF3L27NcqqG9u5YFXtUqFHIpqoVi3IlxUHZ+s
SjN7XcDtLjtZAZG5e91sskOA2dHR8KuvYuEZDPXCrw0M4M8ksXvRIsesmR5KgPgguGU1jdDsYMnY
xMHo9JmRAlvwo23dc7NSH+rlFqgrkQ6TKme0lHb05VfEl3OcaLX1lNqAdCrBPJxD0PZ0Ol54D1r3
Exid5pJWruxaHJtbgZ1gXlYsKPbIGODHwfMXXkhtkli8l2+usDRiAUMtI3P3uhe1ecSwg2cP4w+B
ZR+Y7cCcXwjxpAt2agc8VjNzSwSFWcD4mzsk3bFgKV4CxuDBbYHYOBCZt3PbSHj3BKWsXg5V1bLc
gfQUPzm/7xVwIp+dkNJ1yC1rBbOLXyCYujMRV5AVd6h5ALkiag7CgT0OyMjpXHDc732OKAOKvkVU
L364MLhslNkhkiEGycLwkp9NkGqVs7NuCuz2nOU54pWEf1kQFLdSZqMzqxddIMVBz81swmmdsPbg
aZUZrPlV3H1RW+S6e/OLvN7E8NH1ZkY5h/7J0EehfR1cpIYtPzFwvR4zC/ImvFS5NeF4LjYxzEza
eviFcU8o4E0OddqCyU+aolocX8BV2Vh1A1Xhm6XmHCIi6omg2pGWZD1ZrNUX6OdvidcXVDEccTWe
ZlKPNlashhFyLcKECv07xanYEoSoApz0fCfoajHOhlAr1xe/jkvg5jw26NB1SsyAZWpyjjqbPG2x
8uK52euhuwVA6rM6GGn/hm+bk4AF6nBjoDvvxv6vJGKPZ0UvsmHFLOJue4ATavMDjBRJ2D4GwDaF
OulCW+v5e6ndqeEk3c/SHcSjaRQQRI/EsE63Omy+2FpXm+gGiXxhdCIIHxTikOxuIVj7gyP0I8He
W5dWXVe7NOFSgk14D5DLPIT3UtJT7Y/rRyMPx6UHCmApfBqiXATjX51cT48eU56ye1p4Wc6+4eZM
4lPkS7MBiNZqDKTvrPbOy7EZH7s1JUYcpk6rdzbkS+J8UDQ84fGNfSo14YnVsjYs5LLT5vd4z/y5
59ewO18k5r1SVCOXuBhgzG1Xr6NvywMjyzCSgHwZ/08ml7rc5mpPDGWfRBtxdkQoRHSDwU3Ou+JW
NbUi0cg7NZX/Lc6g56uBbtAmxlc2O6JYT8lHj8t3ESrMqFO9OzN1giJp+9XRSdb4NfbUxPPNIvIQ
vhCMjttrbqtwA8/602ZtIr43DrTHRF8bP2E38MwgPJ0QoDbhU0v00MTBN2VNpi/WXXaDchZKt19Z
C3qvDEnLvcz8FKO8LIXha/y/nDLIHe94ROJRwQEva2d17OrJH+uNv/u29AGF5IiW9T/HNAGCAa8s
Cj8Va/EtUH+V/BOgYo/NYGna6NOefLROjk3Gpjg4kXtnOvle5xJ01RmFKcfyxpTv12vwuTHjtfZW
Hz7jbJiGVgFJoTEdeCDIpj5gkmBIwUO7yOAS3CPHrxOZAFffGvvp6dlUmKQLRrLMkvqApsi6UV1p
wlfTwu+EROkkZvz7J68IXk/H3uaThkwvbkeYVdSpY29W9JjrRAKI8rM904siWmFlbvZJ9QBV/DXv
Qka9E3chojfYpT5IMqGAZq9KVWHJ29oRTUGf387tVAlf3eyU+Dh3SNEkXKqu2bjA0VcPU6smmGqF
vhAdH2yqbgjP8BmRYrekJ+xgK/DIpBe4yQHCRiu4GYyqy0tprmFJlPbI4tywEi9UWWLaDwHgSO8G
6vkSAOtxk4zTFCzBAwNEQthsgdvDEs+0hf8uqBZxdcROGFEIpaWwLyG8yRImV59jGycVNDmhKVzY
unxAbQZ6Z6uiwAFoERrE9DpG9lo39Zm+/iuKViwc5qCZAlNhqZlzvX6mhhP7biz4z9vh5lRjW3d7
kIIbENkQl6t72xK0nSwBktERGjTdjaj4bIzmIag7/Kzuu3p2EUfNc6fghYkV96NV2ElCO+5Jwtjw
4XKjlFe2IR3vEt8UM1oEDTAwOByY6kdeATVsz8E+oSVJlp3J25TtvDdpGOTBxWTIlrIi+ZsJnKGu
izFScAMRBwHBXZxzsk1xGovcX9w7EqHbQZFWh2WfrxXJ0Og2FXCuo3pTE/dXxW4NJVC3pYiRqfd0
vd7lSbxc+HsZz7dEIYrzU95jFnv/ooeYX5AtE2w6+Sow5WhDC05b3sB8PHRsdaRymHCiZTWSlLGn
REAlyb7j3qlTfADXFcWWSTiCnawMxlNgXujzPft9rw2aK74hevSR5XNTxRx0VVOJFBAgndF3LoiB
DPjXpwwy0goF5o850JJA3rUBWvwji/WlehUFpFQYmb59czouU3RrsP1Opf8PYJ7+TvF5R4qKnSyU
P2OQK7MPiEW2FVdztZXQJ8mYmb4PsdWqs/MtblAwqHydwUtShtzTdtpR6S7T9mK+rUy4DDX/Meqh
KAyukFVQNPQD5yOBon4UvJnALAJWfjuS0/Qw4w2+sNbNPlPJVERqbdVJ2m8MwX5eoqw7HkXOXeUD
iMB4soaG5qKmjGANykdIhJ7LZOSwOn7isN8yM5q7qmknERzbgX72xexM0QoJdznmNJrYetVmLT62
PV/g+xWFYqDJDhevoVQc+aELK7XUu0KbPRMXgRjuc6nurkWI9wsNjc12yZduRyZ5agxSZmb0FeZa
4CPvn1KNwPALabL6vmfJitqSIc+WWsnMgDM1aeeUyOrJO/Qp+YpP58CzzXi3CbnCsHh3Qo3KSNS+
192sf+zRmDRui2kwkZfKXhtiqwXLfYI1k4G5BQG4rQm4OpC4nQY5QFOLOMZYF6AD/EJyjF4LD4Ks
Uev0Joy6SwNhdhi1oGcUsT//daiIvaKpN+ZBA0am9Mr1W5mnKdLfBozFrJrO/f0vSaps47bvi4Gp
3D8HZpEecZOwkT9eETeRWYgsqPmHA7gmEhJn7bv7q2oV04kad4v24tYlAB4seXRvrxjnjXgCchzm
CcmlGYzpyliItRq7jTc9hlBVpp36wZSactjHEsAPRaL7Fo9DyXRHLBc0kuCXvDut2hxbNYRpjbdC
nFWFNDy8KH7j726l1Lnrwpq9wk2RKmF9ueL2F1WdtyXqhacukpe2PVeltjl3eI5dmC9klmBjDZax
hZ0K4CEfgmyhKkk4EB8okW0lgtdlOCuIn6uz7ns4VMjrPOa7/5DkeWZzdbYD5OWGoOjKnUqRemAE
QAppvHLv/AKsdWukvF3AQgzoF6uaEPe3oBlIKq196G72tseDlp53D8784RkHFYxc1Us/YF8V3yVu
LklbU/hKHGw0WNI5fKia5VI8dn8HSxX5StHfAE/43zDVTjekjxotaK+iAwr0PVG+ki+zw0g/Oft6
CgD5t/F1bLfRp131tSWFE1EvkUqeeom30NJvwihsm935GYabOgy0qLmrZswONcNvNc6pmEv89xuB
UFJUy9WawsOLlwO+Hns7+N8iNUDa2iPEz4pjKtg1zok2wH8QuUG2EvdUdkUE70+bTL6p3JfxnIJE
oJyEQiIgoWjB9QqIXWQ5QZrGKGis26R5aKPq+1iU7MOXeGWATCciQ1R19Sqm/AWA2XUB2OBh34V9
tQ93nZ7AHMa90CQr4n4qRwlHLnj+INLLmvs7EtT0Ak4AmELEb9RcPyLhle+M+DNeuP9WzBw4xErn
WAtGPEr0BwZBckuKvv4x4cww7Q/R67mSZZuex2ntvdLjYljL/sqbKX2pIROtdTyi0+V0mnzi8baD
myLnG88xw9kYXdEJPq9zAYMA+yO98MvuhRpWvuJvZLtlkqV7KhgcJDKTm83oDrvsnbPEKZ57IcSj
UoFdNbSep3DSstsFmXvUpV0uP3xI3/xlA2/lr/rLyyDuuJYgaHb3tz7k8j9jAhE24wJcWkoPAGWY
wEeyyjryUWGCjcsIN6zwCkQvk2+qrw/kJ85VoZffBqW8V7c7wJyJDgckV9l7vaT4ifKD080WM99N
J+3MBO9hFeJYIlMQXUg7XuKox5zv417dKbFSxy2wgXxa75JS6F51c83IHU/vcFjAWOh1ucQiBGxZ
QsqENXXy9MGJgIpasiaEEooIc4hIRs7+aupap5Ilprga4U+Pgl2rhJ5xShvgxynrBJzzWAb63OiS
eV+NgkNIG0imsjtuR+AW0mU9IwY2VS3ib648vDwOT7qQgxohKlx1kkEZF6xzG/kZ/FyqkTqcCtCI
eT9gCdCFq9IOs5DhyP4AklLRhcDEd9utATrydBVN3cJUpnhrK3jQPaYjsF/kLJS534ftENQzFcRA
RKL+bD4jjcGNalLTSSVWKJoIk4VCSZY7o0ujjbjG/xXAfEVjxpBJBb8FBuKvk3AOkBNXuq6Z/oa/
R554jiiN2+CWhoVlwItyWiL3/HPlZank3F/tP0e5Ee2rPRwb5RqGMcl2sCOmBryVCmBg3mY+THF7
j8doUbxgkB1d/VNKcEnbMewqEgKuJk3CWzyzf6nGti+7zoXphy4szCDM7WxuNzXT1Ti8tPjAirk8
w1379hSnzx9cG/8OJrwOnGzqtuNpIOMewZm2vu1nQwIfWuxHZgiJWOwiz1qqYctL39Vs5EW1t2L6
iwgDULXAxQsm+7EwFpieviVzhwR7fF/OBw75bUwvupy+9jeNLKfrKw2Mt7UTbVSfvAPN92xKRy56
IZMWTyO7G4v7ETo8/nDTM5TztUwjVYtDtJensL1Xq4i4vCph9tT0zzOSiUEKEgkbeEBU+Jv1lg0c
KVAYiDCSNeuLwCcUy7JL+SsU2jRvtI+i0DXijvPkuAVyCwiJU4AtuH7xpgxIKsZMrJNVuoe05Smh
YfPtBdi19/H/A1BR0vD+Qnj0TZlr00taHSJxoWJFJQeBqiYrMmt/57OVyDXpGnCw6ybtQoT1b+EC
mS912BcQdG4H0WhIPcSf2rIfkvoepVM94tLMddUnfqW6wdbWl7quTUVWPX2wTZbtv8uerEonOMMA
ymh5xY9qPK0P0z3R6kjlRNqoINorNt4o2vSD+7MOtSMpTUvQck8I1i84JU2NR9ztqvdFNK+jSG6p
njfZfz3FPbkkfq9qV6fJ8ydKBpiQ7CVNk1ydZBAowZ7SQoGpRlz8KTmBcpIixnSoFTM+REFx1H5b
WgMuHBkAeWwYi2HtSeoVUwUyjmCtA+RYujhMC873iiBwrJgu/i1/JLVfJIq0D1bM4tgI+k+G0eCg
rxmk4VDtbCPwp6hoNWL9g5PeXoOGWvfimHGNENnVTVTXhUV6zaMhgC38hRaAaBR0f72kRuc5npb3
CjkuG7WRTYCBUDVOIcnmKbW6L+yxdtT63NxwdYtEtqlXqSV6USYV4AHfVuD6mWQzdi7uHC4ZbfVg
kPYPBFuuceYn9VcqatnZpY/7n93syYxFHS5FlwaRr2MZ0sJuAh5DfRy3Fnchy77t7f3eCpsKHSzg
Uh/OWrJOJ/sJtWx46O+nOwaMTIlZVQzv+Zoe0uZTsgk4hb2bC5GzbuXdZ4NLj26P4xmJpFqq+1R+
eCYC8FJlC903Lh58cnXmv8oP+3vjim+4Q+/inUnnywEUV9GXhCqzc7miXzj+gihO5Mzs1aAhlG12
MjubV4TMHBvm2CBYydscuWWZqbAAgz56tTisaBsooPrMn7tqRfhvRD4A2YMNtURS6wAC6+27fA7b
lmcOy4EA7n3m3f9t+gW0KQOkTBkBSeo37lj+4K2cIHMeRsiH8KNZQp1JJyOuHkGA4p0E4uZepxbP
D25bcI507Sd9y4lDJ/KmxrWweAy/k+lr6K2F66ET9ecrw0O1UG00uAGriNyBtOSN7AoMmyx4I/qQ
4hcltzSMFcLNsip/k/Ic9SzOJhmXCoFUjZDCWuI5XNeMsGzdnwPdVMU76hudieVjXaix0QzAUNFH
bpWnQAWzKargA0NEnL3NwjTDkqWC3jO4yJQBaBgnOlnvgS2o4od8aQgaFCH8ycpXu25JQ3SQ1eeb
SFQ4o6hB3CYhCgxlcGOK+9zlpK7nrwmka0BkfCGqhsmn+SzGGWdW7EBk+vkOBtTs0GjbG1VdJkTL
v5z2Z8+gkkBRrt/eIiyh/6Q0QlE41JPlsuWIPWGpc7ZxYsHPIBXR5UhEg6H0K7aAILs2vpbEtwMr
FtiqrFC5YVM1ceGoOMFa5gyUnN8Mgc8MHm8pKdj/JCaYfuMPLWPp+YtWjk5EirJWuwp7h+gqXBFb
lBm5wIPDl98fmr78kkWWEHegBXdSmLLNmBXahHLRgXLZ2FADd5qi9SHl2jb20maTHRrGGDNhTxiA
UQNCdP65Iu+773EaLr16LcpZuLa2ExPtIc6Wx6vpfLEW2dDKYHBGm1rDHzfu8CqCVo8uCgx8pBW0
4R+IR7eHp7p5z3oKtFCNFUlgrMVPYiltHJyXgvBV0vAFUoAiYORCkfhbNdNkqOZ2pEcuPHQjSkYM
5l+ca8tpz5yc14GPdiTF/J66IDHlsIwd23R8f305EnimKgQg2nJfdaJHBUdsZDCQan0uRYHLYwVu
iTe8YEMuPARn2nWeppNkPv2NwYwVA7oNzV7AOMyLaYD+ZruE7alk9uXToyp9LzuJqveawpzfXy2A
y7sH4hSsR/w/3gc3bgQZxFCv188WjZjGLnn4zSMbaA1VyFHZm0wouEvbMxW78ww/1SHcDq7M9TVw
kDmfUWhywM+ArZSFsk7IP4F3OnxRLU66YqK0yfQTEfJfQRIq3HPcKpVy4ygIm2s2+Il0wckZqbB7
5QeJQwe/MZA0569N0eMM5AXjX5HXDVNgFA4G5j0FYB1DaZMtXVMI0eDr18iT7lG1VzXGkd5npf9W
0Hi5CPwltdw9QX5+gGFVjPN9geQvsO75X5NCSngqrwnQ0+xfUb0U+EB2YEZwMxBqHOVi4wd5Hbok
DUt4NlHww304uT8Jpt4CNH1AeApRBCzB/Nq8VNnnGeQ7DkfVh8F0GlOUnqS19SL0/F6SuK9KLZUB
lnXjSakqYLWDWy31ZdaU7GkmagsXAR6w/50gxuWQcXFK+QijpeCxZ324UPdnUERhNH6q9EA+k8UP
axP8CtHKXU6JWdtsDGCt/PO/X+eE06YGFTZM8N7DZoYf3tRp9e27CFAU81XgklJ3g8vd9eWKmehZ
uh4F/l1imgKAe0X9B/1xAccRPCzckefU8vaf3vi5fc11IB6Vu66dqPT0Qr7l4512R4SZwvqFzqfT
SV3sSmtsOQcReG0pGUrU1beSd61aBUQkvEzTCnDU07sRJm66MxBbWWOcZtncKz5BjQF+oCvv0AX9
8ySrNcHb5Qo1rBextA2x6pxKk82x+BtwwVfM2RmDWgUl0h/gGhNlDtp5Z5Et4OT4MtAgluG2XXD3
ipFyo3DOW6ZKD5Ji7o1VAGS05RIoeO6kLuxNLNb+oKKfWSYO8TfeLtlZZ47/PCBh7lWnpjrKUQLh
4WSIbq39HRJx2rtJJnokvCG0Je1oSOPug1sRU2ZjeRY4deNuzWdx9Qx0sJfKu2PwD5ya3Qq39eTA
ph324+kxYHhTdh89YoWjX4fPGyXhHtxL3fBl6mmgTm1D08cLo+pQEBbKtn7xgIHpAJzc0XZkW2QH
k4up6DE+g6KXyK/n7lf35nsK0wBqpOzwIoCyuvr7UFdETv2oDGsijQDWJaxZ0kKhZrIn6Cdx+xYF
OUnioODhHHmdFJKRXNeCoPZSSNftRNA4rIRugHlLREHwDz2VX6HrezOFKRf7kCpQunXzfwFPBY1W
0IGcupbtw1lJ7IBUJ3Aq4Rfyajs2o4oui+mFhaHwuFZsq33klUT0x9f4sQYowq53ftpXitHaB704
1oevtQimuSJDWAe63Bh0XjRguXVq/WWWVJM1l8XGvMQdO5cUhL2CYpn1fI/UL8kFCdqvlGDn3MHZ
/v9iccZwQJIRtIaV/9vspzNLqV2JMtcSjNCQp7oqLeWOeK9oQoweNcrcQOVn2koXO/LLRTUpvlSj
7D7ReDXj+cEZKGqiYFDipzNd9AHJxQTPpo59m8Vm4bb3D/+E2emmUwYMeZWDgAWp5kkRwOK1X6Q7
e83U1gTDpRKA87E9PRfbGCCsNap4CRYDTDH5etYEOEZ6/cnDs4lN5vMUUlOri3CsxQDs8vDOsHC2
ZGotGLopFjnAIm1bIMBQZAMYaDPLovkW6z0kSYegmhDemsbRzVHuncTQ6cK5631UjIswEFzYjIR4
61oMCx4zkvlKj0g3pTzUHsDZQlXmyym1bL9elPUY9IsRjM5OHwoI6CWIE5LAwkarCEcwyloPdRgr
KXKD9tJ4InoeDSGDp/vTHFbUhDkVbVXZkvFuUyugNci7dv16CQgybWgLCS8+9ODaDypl96np2bdI
Cx95HcUxkPuo2Mn5HVEdEnznHcr2CKN95ALErhMM+g8RgXLJFbUtHkwuga/O5bPAw//A6DU3nMoN
vOs1kQzWo9aJijvxYnPNrYVYczuM7+KJdAlQ793UKT6OPCJCnc4UPSf81MB+JQSLfxx0dunO+dvV
j5uC50FeyfwYeAzqIOkv2A23t8z8aQBKVUB3LvdB42NEzYQtbZUzPoY2djy4FVzH2OPZM8mrel0z
EeZaTn9hPfeisT0vQF6uahft7HbHOGbQYuoFyVDkqQ1ImAkxvytPrEpsgedw7YGFllRMUQ5rhQv6
7ia+MdKpPfveww3LZfpN8zd9K+MCjytFg9ygIp4B3psbaut+Zqy890DlkLGnoAGE2K4CRszRG/AH
Q57pLsyWvi9WoCYApZspM3eUKJnf4k8WaQIZ0C6vNqbY1Y3RJofQu3e4FGNGnZpiJDUn4VW3pPdQ
YPZpNrtj4Kh969ydqnGWHSNM+5OjjrT/aVJQ5+s2NtuA9Q2uoCOG1jXua9L3NAnVnMUj1tHZ5OBr
LZSbUVc7fyodv07rysaVAvru4aD6d8E3gR5uWnwZLy2rcKWaj+9UfhZcEpCmuyAn5BHGtCW5gCrk
5I54YMfSKXVa2SV5wnByZ6AlBVylELZzAJP74A+3Q/rcHMMyEpqkWo4EdPdOhcIaC9XxSw+8lClM
uyaf+/4xFyU1L9t3z1/nxQWODat1Zm1HnZFKn1dzM4k4yl0f3UYcQE0nv4S9ja98/VC64i5lAj2A
IDB4AQikqyvzGcUZj00ZK1L/r/ergKRJSrrBtVNDm5ZAWI/3gyC9HShIIyUDjR5gXkU9HnCIu80F
lJZDlySzvOiNwtig9DN1jUzAyWBoVepmYqCKGxAu8Ms1T9T/6Vd00EQ+ZxLBgXMdaBHD5RjyDHrV
kU1TZ7ENye9yApOOyORx0hjcPWrjMyyjXgTmvNhMSjGNA/pXK8MIZ50mzZ6Q/TUWnTCqg263dwK/
w89j2KJqGnrIlSRCrm2LQZK7H1+SdmUfebC3Ek93+fym8GkACn+31RE05oQCGymbFT696L8YnRG0
RnQzNJNcQQl4+RHomJZIDxJueZFyKKB2Kx5EU4EcpNmMmyXKbvMSOdyxhROb6gpMzO97R5RVwhC5
FaighlcKA/KYU4nSLIyM/oTCMGRNJyUHz55zXvgKvz6mZarGnwzBHd8FxEziHh947ImJoBpNp5/9
NxHpvJS9wwbQRnFWv2M4pvLajX100vUhR/49iP+Hv7Pwy0VY3kZmgJhWoTxnDLqPSj0ClMaemv1M
V4Hm4a1XI8oy97D1rQZYTQRxm9H1H3tb58X2D/UrvRilhWn+gjRQZYFs8sEXNCN1sGWL+qalphcG
k1a16vQiB0y/DJsnjlkoeytaq7w5Bhl2NQ2tZo7LmsEQZc/YYyFomtArG3MuPFi/tpcCkG2eUBhX
lzpCVUSu8vGaX5oAAY0s/b1sKgROBWIvoA7nzeU6wh5A2ctHp8m3M+vsuCv6Sm7cmVgzXxhewjtM
LcCSWpaRRiN3LlNZi/gusEf2ayNnoLYWXLXfuiY8sfiuZ8TSTdLTirYQFKgf3NAUH8Q9Dw+Cawnz
HsacVfyKexgLh8ePqp4Azcwu15vo1InxemLqZnGyK35M1QdpfN8IJzHbxOba3wM1je6leBSNtO6x
GokefsTuo8gdJ454Pwc9PDgZ8kj8y17iYNkmWeM7EGMO6PdMBB6ppFXYVNAuXtnXh0uq4DFDW6f9
DcRu/ocmORSLKgAVvWV4GjDxrmGf9LPH8jqd+LTNSZRWTnu0Q0E0mNxT5kjAx6R7d+a/xgcNZCUj
Ub60u2B0bjB7lNcaaOA5s3fHo17ZYBkIuRiYDxs0v8pzAnlCvx4SKoP93H7gie3oBSAxeDBdbzmN
lggxDgkqdJaaczj3ax2QEHSCDt1Kesbo4rmPCrL6apdURxTtGFdNN9eqmkeWvaxRamaOEPmZ4bVU
e0V7HdTyZSTGcmHckU+bSFnXKMwhqK79kl02l1hdotpFVHVcP39PDvtW3tyV1tTV7JKfqNjvo0Rk
6XRoIKa7fbKHFBUu3ReafGChb3icWNw/bw2PDD76DOZoGtUqJQm73M0rip80x/U5Ij4vj/ZmlMkQ
btKnPvfVBxqwvrsAhMYORMs6LF4IfT06Box2tvI3emRfDPdmqsx6qgYukbNvJ9Xbh5IgJO7HPoBH
4ZPHx/OlXjA0UrBH92sr2huTALxm42/ldUbl4zvNIlseLEbwceUaNDDRlCWItTGxweqJQPdP7KPd
FzCeHU/alWQa18J7dfyRe7O7W88e3XYuPZe8d4jNL4/UiTlnvKZ+ShtKSMKBYjMTzm9bZoYUvrkf
JcO+0ITC7W4yLQktcESojmIw3TGjQR6oRccouSzC3Gnahq6mzHqGP4IN16Lo+TXLS8NxdwerX6p0
Z/HG3HbWn/Sr5h/wSaOZBFcVDcXPFIhsVRbHD+tQdxHG4BlmZ0XXz6UAluGQjUTfZ/eQsGuZXvpB
8jQlY4sKO2UVXRS8hvXxrYkGzR1kmI0DvmiKaeWcNaGsMvRyLTqmXdhrMLJI72uzeZJvNvJ1yZRI
a9wcYU2VnjAMstHH/ySdptVTG/lg36Y9VBP4fAzclJDgEi+bPmnJQ9ZfaGXQDzMzVSwdGDwKCXg5
+VHbc9/Yx/RmqKeEXcuyizUl/VuhjYfyIH5VoH1ue7k6aUDAJubKqkz4xEOqs/92+3vPCjNnkVoM
zZJIVUemJPeB3Qee4TRS8lLjvmJhrGLnUQzRkAE5lPYCjwzoFATgPRHLsWPSnIBZKTfGlKx1c02k
gDROaWEG7/vkncKuXR3w9BXyqGCfKt4I+ata97G7NHOF7MYkCWZIDCqfwJUCg5LstwDQzhY7lWLJ
j297aEBDt1rn95TRVY0gPTYTvP6WkwPA58lhhg6a+nGqxrIc5Pp8XO2LTeiiBO2JjnHpzUlf9FqB
eevx8gNyzSQQk6lmD4GKZ9t1MhxzFwXcH0yZOHmGuyDXncg9UBbnsi8djuAfU+xHKgoQ6C24tzWW
8oBS17v1ekYuECSoGj0KCcXjeeE+a4MSAW4R3xplWn8VW/7eOvYyOmg3VSDq/6j9ll+7WwC+X6xq
pnfSixT9C9UHQIlGAE/6ssN+afHapd4lSxmT42/jn0eBel7pU+nOWEwcSjEjrM3YqS0lO/BXPu4x
/hfreBfstjXfDmhYDijtDtgnVgMeVvid59zrK+mwT01orLX10O89i0kW84P/V7t5daWqEFMMux6w
o/3rA7lCEUNSqV1dA4bDxY0hV35tQct5FzdjF86U8oq8t8NNYq397WjcMHmUGMtW+8My0vXlKFSM
nmBbqeobmj5RHVfuVb1xdTJyyX8Qwqzv972cckuZqrWsk30BY9CizrDHE0dg9BFvZdEO/A+Pb6CW
z7UPhPnCvpZ4hjX904tR1nbWbyWfZsGac2+B2jgzU1772JB6Z059KSvtc75zdO8co5K7mqWZFyXz
ojMZvh34NfjGw0c3qa13azI3STkZ2TJAFh3BIdxxOI+1SBPLakF0rPCHQ+A5qFRdga4FwUJ06tac
kq2M24RNjk3fsMDwpGlvVstk0rAjO/un710122o1Srtgsm4wd1HtnStfBYbRsle5FL8Yp0/K5ir5
qbS+yxFxnoqXGNpaGcPs0EENdsr1QEp6OQWyFzXYJgCTYh8WszRmNUlUs8UYUSlkbooYpDO8oNDS
/6kRkC9WwtlkXyd8oVhqPbhFKW02X1V96sexVkbiPk/z+jediQSriN5Vo8SYFKg5afCwyI7Lp0mt
M+MCog8D+3zSiZoFPb1ZZqVOSmmQIYEXB4rb9HWwRXH6JA2QtBSUJcl3vO4CrAijlKzydA/JF7LA
Xb9dbgVN0D4SUGxICUxp2rkLyzQuKWjcEWiiHyc2MDoEc+Q2RIRhkFaJjvGiuNuBtk3Yxan+Oa3e
chP6o+Jf965/38ZfbXAyJtukB3KSUDxMO+qGAydu0V5jnKgbN0J7j34u0RKgNmJNifLnBG+I732Y
7cu5iQ6nl7OOI7Sp6ExGGW9/wsPJetUSUv1IJPcwu3FVii6z48pJ6RrcgAAzQ9TeqlrNKxpeMfCY
6ZYp8hDVxN3gfI9J4OFPweYSsyvh751eSQXKXhWQqR3QbaGYeXDDgS1zW+4uMkas8UWclBvXJUup
O5d1Id/+UEXGNN6FhWvhIRNCHweNyWIQ00i3ZAt0IziZpYeHyX8GK6TisvbAYp28GVceJGRKNx9c
ap0kYjKq2rzByYOW5VI9cv9Vy023CMUHzieq5GPolEe0t1d1b095jAR/MEhthXKruOkItnNwPz85
Q0OMQ5sr9MTsKcjzn5+wb0eEBFFhZw51iRvS1Sr+na2hdw41hdQh+skwKvddOiZJKFej4xVf/U3I
78B/dVrAXgVFovlCbnF6Wt46V9Ov1E3yMH7vElb1VJobTIKK2nTqc6yrOPn2U4L28F5wVjgIe4ny
ra7ixr98O3JWeO6vix0dp63I8jYw+wKRYrvTvHIEVcRiIEAReAx4c4gcIJ+iJMEQo1jF6nuNXTMX
SZzT1R3WxVRf95o1WOwbj14qqE8vJH00dlh9O0UQxtYw3Td41kEm7SG6OV7RDGu3d65sTLaxvkEr
q4rvcJWUa1RUwEr2VeGgN9+fLZnWFXCBHpOIJz/+YBMP5x/oGzCNhZWa9OKpZA6RmqqG+fo5jyFn
goxibRHnsVtgH2MzaSG6sRyxJ90JjwXPp5Oc0i83Cst+xs5148ZEGcRAQdjn96AJYlAOzynkcQTL
rNq6Mo8hkDR7DptcV/u+SV1CxC78P0sBllFl9g2bPvJSGZyqTUWpLsnn2dMUFz4bGBqwBDTyRqw+
MLUIX2270Fm2gO+ilhsAlUGNC1EjTYiD/Azo5ao6OS0c5u5SLuAitWiI0mJ4Ty2/X9t8CNbdds0q
cNMdocoSN9jTaKEOYOEVOIKiKghHUqBOHD6e5/XS9CxxQFi+XmzexbNMvo+zlsW9W6vmWtB1/HxW
5mONGqSH5AoID/2slmEXLBEGeJSBxw5RUxrciwgv++5fQUwzM9X4CBlwrqU7X/wGL5EvQGy76yho
h6PMAbeMAA/GFwIwGNbwBumHoB9rJe3W2m0Wv9Jsr2oWtZpetny/y89Pe+C5mnGg6MZ+dHg8eYw6
9gsr54OU4OCjLvk4Fq7E+iQG3K44a2xlY3Mqeg4TnPhmx8Ce78J/wpc2zPIUz5Ok16pHUp7zs8iI
nykgQpaiZtYuS1/gaA+2XnC2PWaKIn6jPZszNRAypE/DvKXrpOVt7sKy+iy/YJss6pmef2rFLmdl
DFn36WAUetbSzcpQy3VJswytZ9lv9VlSChf5ZD/tLvE8hugHfLLvJtKzrFC7qvaMwgrQ1ktElFUo
wmlSWKs9VDCjs36YsmP4/dOoAtrTNUmHMRzQeNlhMEF/g2g4ViRBYxOZdVW3FIkbtZhrhtEXVkix
7EwSzjioZG/o3ZltimVk+SOEunZdAuOsXBCp6zQiz2j4+rpDfUd1WxsxOUQlBArUwj1r7ouhYcZh
MOOPK6vxRTSveZGY0iSNXDwSgGMQe3kMOX53VpttTFrs5CljoRy6r/f0ql6gtiY7+PkcQkrV47/H
p0+aN3DtjT085wYxSFmPLt9SJwM3vD9PXobId+3elc9P1yDU9UOOx+vWIoPO+Ml7KGezB5ltdVHX
REAbZnkamRcdlSCw+29j7cMcI2sTLPLiljFlS/6sz+mTMTrUaTFZtWgetkwNtiSrQu9LMrhWgv8D
wdvWorWdD4TGEMfr4Yk4aZdIpkOLqf4tmw2nNKMuMftZOArqAdHRBtbY+YcMid2l8Yk/Bzkdt6tg
yXbMXr9CdIvx2PEEoCkLcOoAIqw132z8N2cR2ccYckNp/1WgT6wLVpHvY1LGtOWXq2hCcRgOcG4R
yeUTXvMyKT2Gd5IJdSM7jRVZcwKh1SMZ4+C6Qm/w+6dE02odc1p3Pk3gXdYlZE8biVXJuHYqsFEq
ENhH7uALZLpqsW48b1qQLW9x1AyWlV1a4a1nwrvZWfdO4ypleuj0aNdAri34CpT4SBkJCSshO7r4
0fWE2jOHnYcmchbsUky8FtUPTWjopOJUDSLajBifnC40tTlzbFd60OSSBVzmL0S5h7MC/NaTUDcH
aZ013zaSuffJ4iIPvRR0DUFzTxgmQNGnRkTGDwd6rTNdg86f3ZowoEAaeww2i5g1soTHgNfRyTmP
YP7n0ivcdVeAwOD5Dl/6ITdtXZhWJzO6U2xXG04N3Bb4YPvnM6re/L0NfwdYrV/nzG2+15nYdYyu
k2oB7Ep5PIGBejPgnJzuZcPW4YzrZhDc0yH7mPX8nRKhJAKLjYGLdrYKrWTSYZ6JDTEPuzN36ynK
EkPNk7lRu0zVR3jJQVKzow+NRw5x0qnBQ2CzUDT65oOJy445nytgTxIGA0VFbrHnhqu6Dg5usImv
4tbq8TduQMEezcETrxTVuIQsPM1R8adVX+iqEsF4fg4LnRMJdy9Jl5FRafw3vrrYJ3wJxnsUYeuH
KlgGozY6C6B5xIDrBgA4YFLrQ9I1TSzsOMYT55L3BhLWGAgTLbboUKm/jG1K7FYlwhZx0shfyRf0
IePKVpCaqC+hu6Kx2zXfp4ceHjoit/YriTuu4tHjbwaGZjSMbY28LYUC18grF8dq13yzqDQ1rer8
WGgBToAI2TlejYqhYbQDbVlY4fuvp2NtXwgpdyYEd0CsXHK7A222Yf+9/H/OxtjdvKDFWzii8e81
hy1zxeykQNBhn4o7P6ccgFp12DZPOnQLCasGxJVfSBaUn/F+5OLCrzIkXeVSzzYX74FMS8677dQ/
XGJwXL15YvJpFevwMzt7ERvChA64BzTsYpJmqMWmtshbfta+vQPKEZvinYzXe5zHlc1mcSo2A4Ub
Cl0j6MW4hZqP2BwOgW3/Dh3Bb/Io7eiUvWvsdOIhdp49p7nFO0OZW77wj/r1Z+9sYUZO+hanertZ
no6ki3juRIVnfv0cgaHa55IsYHx0RunJoUaFItlM0LuMsr20reGwWt1QAjymWOp7JSo2mpWcro1P
o2UpI/UbxwYxcE/OS8YHDJZXaeIQOUzeQxZv4kofTZOeyX5alpRsREdfnYzkyz4qOzgL/IfUG9Yc
fBzIJiUIqeaseZQVkp729ATMlDqWq0kBUE3L8Bi7RRe5Uc4YbF7WJplNPr+OkPXJQduyAr84EwVg
c6Oe6u0KId2mStF33RPgLb3L37c+eJmrwARvLOduUMPezRSyRZwCUALAOGEQ7Lu8TH0ryGPPzQqX
fkceZlsG/8uS/qE4nh75KtkJ2fenS3QNo9jhMHNMY8R+haSY5o71EWvpCGdwgiUrmZOTph/aYBdB
/po27SM2Ob3ibteW+cjtYa5+BtA9n7uKzW5Xar2DHZRIulcxjYGKJ2HoyQ5jba6xiPchYTPOnBxA
MFq2jXBs4KhTTmK+XMolAYfXg2RMtEJnLhqTjqR7UPiF5HJMzGJ+SwC1+mnOyp6Elz6zDwKcfCON
5HP6S1FigqEdHrK0I6UEC0lgwejSaxy7SwJavDbk8bUoqiDLzX5/X7ot+w/+vYI0BdkVoQbNUlC9
vaMGphiz+ZnljsmQVdz+AhXG8JsHKl8diAXhYxZGineUhi+7aHT5mgvqGkOAi8gcm+uS8+S54Os/
5dMRUwKQ0tD6XAUhQej9w+55yFGyAhobr/R//vInbpoEbF3I03/eTFoRaBoFZMOo34wT51xebPw2
C7upNdIjjRsekuH7dK8q+SU+U7ZM1BXty6lKPL8+HakYoWZPSzyo7zWShzP4/BvY8B0bMwhTf6fV
ylk2y76jZ90+SkI/0th7PqRvmaQAedxE8TrysvKO2qGhxzONID2t6QrErkQufNRGKNqxXNAVGccR
naYtAEq5WNTWHpMnugpcRqb4ihJvPuemDet8VHi72Q2TE9UavXvYxpEcXcDT1ot3GXGIHxcvVlld
JVjBK+oRjXYcM5juNmKaTT8RUa+UVTsxE+i9TNALgosrHSMb99l4rVAcxzG6m0WOHuJOjzBlJtNB
BpZJG1+KjdM85spRDPrl523hhfd+ZvLYObrd4VdXb1pGSuFG1/inFh2gypOl6COdKNditlMg6cpC
cKbMvf4C/G9RXaGkuOzK8o9Cqh9Z6uKDhRohz7nvkeCV8DtU5jLZo8vfkpspiMm9ccwvRwx7QzUW
oI+FZwBd5R5/bzbrxFV7xb8k5eFGLHx3cS0BPqhaPJvLz5TJh+UNittCAXnjprSdk+U4cnKRqAmM
ReqM4PaSFVpSY5aGLrkm1yMlBPyr+Fxe5Wi8ADMsj2eg8tGdCa/LfBXU8NLm5/THqGpJqVQ8w7s8
mp8GYpc1AsYf4a6HHnQIYRJeisW4lHQK0FN2lFoa6qOtv3zT94GHAkhKRGyayNLiinnJH0Rzs0pB
1ClAYt3ZSxZ3CPuL8A0ZnfNJ+XqM61wdA9B+I2LCZFkR/iAc6F5HQZ41PZ+us08w3iiE9F9J5/nl
4E5pVM5wbUPuVtIs6NhJPhsZyLO/UHSJA89hv7IQw/kpBatkoNSMJqQFEslZRNqAQCIyi8Qsc8Tu
Xn9xBxaExw47rPBD2S7lQcz5yq+E+0sJUt7XlpTIZu5NPR/DdtWoqTK1lfp8Iylalr+I5Hnu2fB5
jOyqXr3eymhoSukej3bbax8dR8GYtEqsrvApMAXQlaESYm0vgPE8u190gDgKBo71w2B2Xh3+Idt7
XhpVFhbyy10M6xqZkFsffqdcb+JZj/pN3/ke2AHRxA26FtZxeQr0iL6Xy7qNZZ5ilaNxSHzSGuG+
zOWvzoksKMdQmkJ5NrL0HnGbnlNHNyo533w8/JmE5yU8XgNsQ44upq5oe/K1v7JZ011gfUK/qCE4
G9tT4MD6qcQNE5Ys8QNyywsUoPCfbJhdUc0MbJTpswkB0/oLQUi/o6+jn1cssi0R3P/w194OzHXG
k38VwBJ1OFHYlpVJYOTBgWDAtyxuX8zBL4ME6qFEJzXKZcFJxGZv3e8AFFnkFI7r1mFyvc8g/Fx3
xdhjCW28j6C6POm+GXJ9ZcqS4DkBMFZLUabvZkz55yKNDA1qb8mB21kKLb/5KQsK+FFxmWAXr6et
JXDfv3p/oiFBRugBimvw3dClVT+p1Ahy3dlogzuuL6YM6UaB6CaWxQ8QC0djYVK2hqFgr+F6++Jb
GVK+fH5EkbFmUILUrHUz/idPfF45is/HbuN0ClKVqhPDUMB+8XBCGErlZz+lyeF/ZHc84VDTTK0z
X/xDVfiJbtonFzZcbQAfGyYQfWW0aKJrNTrvJSOZy3DH8KjSqQ4XRfYGNACZgqUfHrKW+0n541zy
hwFDuL65NLjnXyBWZGFcmsKoLUzg7y0XQgpBIXpEEaHRna0rD3/vTxz6o80xLtp3z/f43O9aBSmn
pTNu6Q6vEiu1C7MKKN8GnGI9jSJk92fUFDmDp+ZH3qkfZi+1UPjpGCUmwAoPJKnWAw63G7kTCBRe
s/HNtmocNeuMM3mnaTOftX6/nUGtQpbo828IWQN1uhcHZIOYGA/6FOQ3cAAvVDo+5zq819gI6igH
XC/NTr/C+sU5ZB73DK2+63qwF7IPvaZlFSA3TnizM8Yk3ugdprEd+WPBe+JGUeTeT39WC6RvZ1F0
Ysi/egZAOah2Ih/5CEJbVGDtZycysjf1HbBBmGJhOYMqykIkLazOlASqz7q8B7lCQ6K2iOwPGK2N
+7FW5VEEAZcC/Bx24z8+KIos01aZ/IURqwsaV1Suil1yIu91FgqgfXbZLUaLQI1qsaoaJrmCqlRU
eTZ0f53toQiKVDZuChzrFwQUrbLtkANh2kZxG40iEaLDSizkg5Czhlg6sdtuSUSX1I4K8uy8uBqM
aW0Q5y4EVDbcJVobNiozrJxJu4QIxoGoa1XgFsRKdVbryOSa/cQnwaNWIonCLdwzvGCf0AoJVTi5
j4m1jUj4rFT2wvlF7kBLv4UE71SqoaIU9DMCn4b73RWA+3WI9GNPcoDkL4rVPFC++XNq+IMo/4Zs
kzVVFo3dI5UeCjhHrFi1Asc1Lq+LnY+HICV8x5CJ1cpS4g04UdVthO8VQVn/1xwvDeUtaS+K85k+
IntKvs/gMR1ZBZHP5ogqXxov0o9x5suKG1wKHlbDbipmqCNaqJ8soRQcOvSCzH6EtikqJFhqVTuK
7xcTGtF4e3tOwbcFEHZt21/3oQLteRJgx3ehFKhg67pbex4QORz872sOrKdalwJEt+JjV1TvFghM
pb3oGyenRybm5OXNUBmSQquMMgpC9n8nKtHVrtJSvOlt2z3fG6ZJ2rxriwDhQq7bDe4U8nMIK+KP
iXm9Esq2BmZK/d0PU17jsA8WmPio+qIOHiH4rKCePWdwMjaR6uePYmvM3J+XFmI8rbHfgA1Luwy4
w+qQFJYCDONp3A3+Gi7OGbE1zeGhiXdD/SvUfx6euU7HeutbCFWzkqxaX9VXnHiBo0rzMt3PlY2Z
qiuk3/+k8AmGqAoigaFaquoSl3kImA6bmMfT36rCsyRPtDBKZmGAhdfIfC+yqp8/bg2OjhXMxAFJ
KZhS2QHDVznk+Ex6y0SBDRVORR1iMKkfp+kNLOe/9C07CR1yVobI2u/XalYSgx6fY4kjc0D9JDWg
zV6uDp1f4Ay8hwIUUADS504IUOs8fYMSb5kEuvVut9Ho1mPsiqA+cMfgHoP2UahNXmV8ou/KV5DT
eEVN9StspdT4PCkYDxdjzyTh5DANmI/atcqHu/vz/uqy8XgFRF67nsz8LMMgUnC+m1wKbnyDQ/AE
lBO8+uZHpgXeyYY7brSPlmLhJ86LPiDGs7Gt5DF32ME70Lv4fyjnvTvZT2rSNIN7C0RJB4Ij/vII
+ZZNpfHHDNtANwHC3/b7p3EAVaQrpBCkNQhAMnkkzG/CIf8HG0dIhQHcUpNT9xWVS9xM17EcTAiQ
XnbMRcsWjSv4HzYkCZsqPCgzuYbtt5BnKsEZBoSevXccjx+KzJw7fRrM4Dp1cSnsTxeFX9MvvOZk
5aVmp2DHgFbN9q983ORSjJ3ZulqkyXCpMMSJBQy03DrPVZoOy6aOJlRBJycHhBjrZbv+6j9XKNhr
dpSOGfpqQ5iP3b0phDEu/DPljKNYFJQTr/57B++b+D5u7jUoI/NzX+/lGObRLZlGr/MCeUS7Fyvh
is786Q93TzRp/BeIJv8GftKR7r3VQci+wGnO6Cn2QGvrcdDLTDeAMipSlsdKWVERfGOJ2cLDpaWX
q4yBzsbbqOrAwXo7b5vKsHFBGnn5n3ILnNrimqcolBHUTnlsw31KkmOmdDvshU2mCFqRMVabfjUw
HHhboVSdPFW9uWuNUYGeZZ4kj3I51Bj8n4fpXC/stsap/7ODjzXPR8LVWsgTNWsdiX9u4Dft30KJ
iIAXlvgP5SdD+oTGtnVhG42e/6ZiO/vmx0M942jbOomMJa8VrAzF4GyYmUArWoXmgEznDGyVWZr0
Dsc2ij/BzInAAXd++cGm53MeJrAlVr0Ol+vdKkF3Iz157PFIYEwdWEBylWkcMEkGX3M2rv0hqFvB
q/RdCX9pwm3H2uOYGaU3XA9xtCYZUcTZuryQeWyNTBl1+J8F4K6ygk0ON5sT0yTNhUNhc4eyX0SG
nwKMOw03OMsATfkEknqMihhbo3iaes9Y7l9XR4+FgvSDfkZAZPOW4ulhDBfuQgwanqrXq4Ogt1Ov
wH9m0HV5+IAxJITimt7aUEbZMKUQ7/cH70ChPX6/nIIGLSehhaELkR+fMnfK9D28kzxJvZPHqWZm
Z571sxeTlLiwY81ZOqEfzJnGmsmBG1hWdI7fy0EgmBO+cyVYTIbbDoa+LGCnDocmqjDAVDT1qOZ6
GqpgnKSXeB/tvqFADhgiVTgsNgZfdnYLuOjF1KBqUB7WHUPauH4Ku014vSDekwAsCFERCuDqTlAP
3Gr2nIu1x30ggHBeS0hssBLbBdNwlPDzYiEcohncoSt2Jz3jti0m89VuhM+CR+C0NwuztutciP+y
tc4qGMnAjx8Lt3zAFmlY7xEyAMRakusgePt48I1JW3V1y6WJsbkDDL9zkbzqKGirvbF+7AzU1lDw
lylpFVOJn0kMnmdl8YB1ZwI0zXxpsmJIanD5R0tCMvlFSp68ifcaXCbJzPnurIOTs6YjesoX9OKa
yttoZc6fmpi8Y5rMe/6v0X5IzeDMpDuKcw2Vzcz//rWbczpW83oT+7VyupdQ4yi9otOGGqPLTnPK
v87nG/2lmW9KlO8NpH8/XKULuRRilfsnG6522Oz17OdKBkCRiCdu8k1EX6E7GM0em4AX7OBmka48
2RrH5WUTIKnTMorEr6xjgJuZr/8/dS7l7J3uSWbs17oBY39zvAoVbt9XeG40dpJC/2R2pIp+lkYg
kkUXpkVCY2VvJ6IgDUa8t8yw3O/n5Fdu1d4bDdboVngYxQuz2NQqb+/wJeA+Uo5dLoOfMLBl7Gb1
8KcHHG2KndM+7zJJQZAEhkSRbeD4TML+ADsSpGkp8HwaRovQVYiXwjZ0ds85XXCjJEyDL6X6Y6Hw
ErI5qFYfKINLa19WVEFiw1egXIx2yuugOl8asxkrKOf6cXpYmI2b9gqiIX7OisiKmLsXm8x67hd7
BiUrNTzj5FswFX4Ca7JCt+tUu6GmvQMWCD9Pz/82yWzRY4Z6yavo+xqsYBxQvoSvq2yptKxSbnPS
5SYhsy3pSM62kUqmfDekeg0IRd9dc5/8KSld2L3jMSuZkIOgCAjHo3JGb1i1q5JRaPtd36KWjkUy
vSxussycF23oBL02+/MeGC0iRZZP6zzRsey3DUHWrCMwJ6txWPzH/ETz/xdc2SQAldadbHfOuJNG
kkJVrvY0i1qKLjSZr7XdIoLBJP6ctfXM/0TLwjX0Pa3KovPy7jjgOKYpSDpuWViteoJorhXXgCuC
jusW5u0XxtJNUjF4jRq5YisqamWhqaknRcNxSm7ena+Z0v5RnkGa9s3OWJ5SJCIpKqE9RXmkrQqG
7DYRwpx8V/wtF4i76GpUUfzedf6qz6U2zIbBLgztlvPEG7z3S164p20Jb8JB/vzAO50DhxXSiJW5
mupGrMa4GM4h4Z2J14AgruIr279b5wnDj88zmbUxvDi37xLS6c9efceHaMGUlVl3e5vnLhaG/WJ0
mQIWeladiKgUXhQOPdJrkNSzSkshJEThEeUPzVByTvvZUhb9X9l6c3zjIfLOALCIXyJKpA0bBCX6
1cDXrCbnKlAR/rdCFOHgzgK5zBPna51jAj/bQqWHPBx8TouVck/ryCvqppQUWBXl5FR2DK1L+pQc
X+E0TBJkzvxsorYSWQJTAWFlVf4PsdJUSVv37au7IJMlEeBkL6+XO+EcJ35dC333wUG8WJnv7lBb
FbFld4rz6aGYJ20nEon4WCq6KiphGh2uL4y4t6Sn6oqlfsLvJhczTrqZwAk288I6zXzx16DtCrFs
PqoaWRLBJkFIKl5Efm6q5ySSVPRlnLsWAp5ZtEV/+dcAYdE7x6L3ZeD7UcZUYAtECaB2Yg1F9vrY
Y3zFL3dm0Od6LubOjEEbmA/BnwzDG6fvUXOJ/eLBkioQgPI81Avoj2KZcrh85ORYNG7+qng/rcxb
pHQmBhTm1b/9CcbxTEGQHhtCQFyNAPMmkJgoUp+xFmk85KVMA81bVe8OBBnF9EDK5gXn/EYDtbdD
T9oxcOBq0uOQyl8xauAwsqGjvVsWj9C8RVmwjhIVj9RGC36DrKHvfdgkysVIGdcNHsE0spDaXhe5
VwMAj/1WUOAFDAaC0LrZftUF7RKWrm3SmAPTU+yKlC0MHdcuZmBNGEkmzKitr5do1jo9mI0egWSQ
6MbF5tNwbdE20seWlHC/RARJyQqsR15FFaxDSRCs3+6JY6HncRwB0TLJrE2QMxfmY+o2FLPOpoL5
RPego45ptzRtnVTGdavh2ViyC0nv7A6i25j+CtOthk3USMqqeezU1JqqPkNohqK+fS02Mk6j0d1M
lWzjpE/nS7AO/fKqsjhh5QAfFMWsvpRZMNsUUloKUTdGhYo83RfFOTrUBL7VadeJ/JZC7lun5Vfg
BDmDSbubAsIQDRue3ZxIe37KwD+yGRox25gyzbx+1lIVKFBXKhNSzDmipyY/5p+GYH+nZqYLuzHf
OWw74xXDpe89MOImhbKMH07OMtJlF2UKU1ejREwBna6bhnm8Yea/KIYPJPW/zY4fn5B5g9j672VB
hDcM64b3/iXen1wWsdXtkgikPDed8JnmiTfAr2YOOUU9fyvrrtphKkx7xxhE5ESer6/49BORpRYk
Om0YhCgDAXIlE+2Kg/KKXgCHsUNHBb36MxCJFEjy+th75zcOPG5153HJF3LoDj6q76X2VLfhow0E
4ES2K63UJMQToebxNqTsdBDt5EfbyulWDpWwaY4e9clzL8bCMtd/8xNSQwxIgv/hogzIOlnfvqsa
FyR1b61j9AdLbORTn70J+My7hvNhPRZl5kliHSwhkJtl5UjQie0nNRJVnufTaAFtmw3RMcB0fDKE
Vag9fAg3eWbq7uBZ7WY3yRy1WYnsoSlnS7F+HEcVqTEs+Oi2QmsC4mgSNvENlHEFZiHP2sWzpwZt
E6Tm4KnijRb7q1OJeznk7gXNu4cq7FQSiQaJs/s8KnTiO+yMOzXXsYVFMABJqsMaL8r/Hpoj4x3L
GC8MeLbhLH7UCPHUXUR9GxICF+AizQdpBaL94JQCfr8h9p0PW5riAtytZ0T38ZLsDP1h+prmAclg
BncgMHpBwe/8zJMug1JQNJ/BcEIqKxrHjfd+ZybggNKnVAeKevJwy6gxzjMj5dhE/QSaZXl1vY2X
wcmfe48BV7k7oQZp/fYKW0que8y+3CKGQIUU2+2u3CX+LgZuf05Nq6sTHozRMzIKtZArVTgAKdEm
IWWsoQ5aYPQjGBt39j6qfcP13izKnKVbnp/pVigj+YD8fMAyApFerUntU/xQjahXqXyLusoMpTyN
NZgJzj4dyxpKTIP6gWakQojgEHxcKOj5c8iSnBQs1/Aj8hY8401lz0KW5qae6zA+3Vk/mR/SiksR
dqKZq2OecNnL1+nTHwvHU0Cdz6qslmi0KOMhzuPfGL4PYxp0QUVjHqXj3CV64gP8Nd1/9AkEcPOu
JvFxVB3taAumFqPEcvjgbWXOEgwmAIczUwqo3Q3GiwAFODYBmsbYF6SFu/BPO2LTYvwwXEVV08KE
VPaS9RpVpZ+bLo/kBTac3pIRhpq9jJio4lg0+lxtSqsdPwPnJ3jADYWlVZ8FCjx/7RgrZdVeKxEG
iBXMbTE/Ks7JpvzkLJvBcvEZNKfRKLeauMX59FjpHKwrCJEydkGiR+WrCYpDqUIbwdOinlmdzCac
nJY+KuW3orDNQ7EGbVqz6SXT7SQJ9/1UikhF+luILut4Ym1Syt3c8UPS35EPeCIIsKIog1z1OSvu
cKV9k7Vdk0DYhhBLAgtZAQWVWoQmswONxSYrfvuL0VkudFBtCIWXaQ74HB+CYtVqwZTeAY3bqVcZ
09hmgS/jgQuwy9UGm+JJRGd9wBlB5+sdV84v6YKvkLZdoQFe+kxDiVo3hIERT9XncLJdhZQj0+/I
M/ViKkqmfJH1DMfp7yQL7yYBvBmjbEOXhJy8tkbEpKkoPWvhW3tT3E3o+hcK6XvQGv3Z9e1SYM+0
9Gtxf4iGH+c1S8OzXSIFh7p5bs2DrncVNGTfBPztaC4UvZQW/2hG7S4Iq4zoxxQpGELmd1YUlUzZ
25bIcSJ8HAxHWW+R9HlSqfc4l00Nl1Duq9wXtwppXYHUjHYffZivJ2I2sDYQmHEsgSteLYn/KWjd
rWFsMtCtEO7shnWiFo+JmLRhH3msoS3ykAK+g3537MrcCeoshJk/oo3vcwML+LBPWiNjtEghylfA
GMYTyMWCe1/UUggoUjw93Bj3ASiBW2OCQd8A9Zwa6MfeyGFki31YkE02vbj9vb+6XHzvUWFt2cCt
xciVvYcPtgPKc07LZ5udflXBOXAPElyNIfoOIQTB7lnB94PWkE1Gbf6tjfBOIhdOLFSBzvN3/N6J
qX89O2LBdYeSAni6jdrPT0iejAbXri050JigHlKKoqTbYUhh5Ofj72VvNRZhdEL6LHML1euk67jc
eMXyWFo+6f71vzlucSgjizArDgGLzTW405WQgm2q6i/wfgXewKcTrLxXrGY2YS8ZyqDA1P/8Vxcu
m100bUoHo3dpo2Zvuq4Nveq0aiDPXhdQrtxJPYscRndxZngsL20e4bTDFO3AMYg7a1cG6ef10pNm
8b0Cgu2Ud6l7ZwO+Gs85eqPmAa7oq0VCZLtrLGti1QDWGnN5HiJAY1MEzDoUAJresKjWEBrUshZC
ZgXPGo8nFLbytj718xWDb+AwC24OpVk4/QpcHWADdAYdOU0N5DLOQFSJmrUbDl+kwYRCoKCgu/SP
/BsFs8F1pisonjKms8STLDmHgiGC/1nfTBa15XE/pSPQLJGFkJk3mciZHxukqk0xhR3AeeInXuOc
SIGZmnrz0r6sZgOm241ibRQgOUs0iFYmMS81RrDk+8G4ldU2dHg5Dhyqt8lW2l9/rnM4X/hTvlcR
0CqLoDK/3dENQWoqOiekBFj7Tp/QjKzSVQN9sWc5x+CQm+RKt6mGJ7O7YvjCJgKjeQf3y/BHFeHq
E0QUrtvQmbdowJNfxUv1IggzZsDWhwL7hpL1mXmZd65kQwKEANal5H5KD6eyw1BM73bcKmthZ5tt
eWWTSyNfOnXf3xeigScOylR16a4QRPa7zLqkZTn0srCxyh2Zr1bncyeecgyQd2aR9q8qGPK/rRmN
+RDZ34hIILg+CBHpC9AXS9FzdxzeVpVjEWEnQ50CzULL7p28/QgOOXDdem6I0JvxSMVDKP3Cm/tm
g6t2SFqhQHmbM786B63AcEkV2uNSsex6i5ygr4I5Rwjp5s+KIdcGOzU973netD196KeHXWUleOfd
cLsbjFF1NP0I1DIm+WOZUq4ubv3x9/0/BZEjhlxDXqglrD+qgDzsa3Xvpfw0JDAPm0Ga8tB4c2oO
xy0aVEMlWtyrwDFTRt757xrrReTTR5A0R5qfLggveUSGRLbwCdgu2+Pw04yAoc03q9f8tgvnbi9f
ujP2soeJa8batSVZO6q6/qZzQqGM1RG5OyIKbaBHj0AS/Oa1rMmuuoOmmlFXzPBsrWbuiXUeYerD
Ev6VUrE813LPqlw6IkzzE8q2H/3e4gMA6qBETCzpMmRgjotoRmlZjeh5ld+cMr+mI09kWXmLdJAK
PjTjGDe1KMUoNGdGB2gyBrSIdmiMWbbJPuSGRG/M2uyslfqChXHzxeTV3z36+2Mmnxx/9+TNGIFt
MSwLH0TAt0Q6Kk5wxXoA8afomBCUex2CrKNuUfaLW2kRL181VkBPdAJIVykrMuYI3iPashj7vLIS
GERTSuaRx0Nhr4oPaxSKxHtaBY7XbTrN+f0tItH4AdAkVYv9WIgUGdziduaSeAZTEEqzocOOY5g1
SlZXWz8k0QkaIPp3zeEdw74v9sfv/+ZY1TO/ziKice3NugW5rXx6WFBkMLBC/2fFh2VQbL4rYMcc
0YwTDf9b7ycVEdH09W0W51lq3GIJiEjQujfxTTAhyezX7sFcUoIbiZb3gZBRZfEC5+Y0pYADP9ob
BNEgpHLx+eSbwyaccemhz1c6bq9P2xJ5VwleyAsKhOUNw513NgnQ4kNwSuuPBf2jfpR6CBc27nqt
xSZ1f7c4hAM8aYATwtiTfTNmcYozudTkvfqT9+7m6o0z8oTKfYx5aTSfxzEnBML3apnEyOGskPxa
oDnO/Zfc8uT2274zcKofYlRXYGuytbCwge+7eyGkvT4td+c2oWt4Rh8NfxLLDTLlekdaE+GgGYI1
6bLfaeWiMEiaEHz9ZdV9RIx9oLaR/wfkaIEKlzdwWnSFuqPvl3qUH7lC9iKPUnxra5QasKGTxVT2
2NtRt90LYHhQ4dKl7wHj/WO/v/qE64tOBEutIPxnBplwythEEV0WxINzuLxJlw1/si/mZsDB20Ca
5UgeAAvmJWCvOEluM5h2jen1kBPF8E6Um7qwBDXqy22SaB1kPuBTvNPFHCJTxDHTaXmBhwGwGds5
/DNOsCZC8G3Y2v8JJXG7gkZcVKj2ROsegYVj2mRv/QCBZSIzhJPAW3IENXGotfbInajkvRa3p05g
dyuGNReh+lQ+3veZpKpa+4ucjjrjEMhVf6BUXkWimABvx/LvBCR5NqoIkmHk7Az7sFzOBYzVyVGA
xqkng4J0HOhwHt/kpzLrQzEc7xDHPTQO4tqNXlTkhDRwRp04EMG5l/6fpOv7/qXIOYd6lIJuB/fn
BLTnCVVhaKDlmlckBWxTPmmTW2SnzAirkeAL9kKU/V4nMuXSCiMaOKjxW8zebKKW3XgwXI2Nh+ad
rprrlLAOXa2rkKdmm7Fbnwdpw+DClvPjYYlbwC6fbWVOHNYX40Y7GRe4HJUmvVmbL9at97dAlntO
NYTIyZi4nqSJ8frA+LsQCMYwgLWTO8rpwWakFWztb3JlEltu6qUeE7grFf5Z2F41D3AueojgtdsY
uKIpJqjuYOt5pNJWF//Yottso6pUzmiI5wvB6u4ducUgrBZQrKEpQxFky9EyPsSnOl70dzGC75mb
DgVZEbGjGAVtqlSsMjtAj55JCfp356kDa/QiKcRU708lHpt4kCXMt6oP9Jgoj2ZoENr6z+UfgDtc
Xe+9u8pB+hxOILBPYdgRj6cVKe4Yayzez3L+p+KVJ1ntKU8d87c6nR4eWGTow337t1M2WQpsSVwj
2sKhLftcwhTv1isM6l4I8kc2fCmZxNTRBEsoDkFxP44WQZclVhlPeh4mriegK7PyY8ThBMwti2+q
ReKdZOL93Wt+Jef7t+LbWDvxTk3FIc3NBsuMz4cA2KGdYS2a9HIlZX0tbUJ13wBX2RvKIEu/2lWm
rNAaGrYE5KgloXkpU7b+kiQgA8jseUUpAvbYhCtc7nTNL2p6og4zEldaGu5rzJFRnllris6APn0A
HTpbri2ESQIc/WcMw2H9Eu8qk1OYWMYaplU9IoPB0u3ISVZTjYlRHtZYJg6EUt+UtgwAxmdPwZkS
JMIai/k2RtY0qFoyPInOyvzPd+MDnz8A8tx3yj20Fs+KL6Ob920G43FOkm+FKTppDx1gCtc4D61S
W/WkFQ1yVgbfwKPt7uOMTEv62h968VTB+Acu7D90//9Y9JOZwjjXf28xtdL9ygMTQHtK8YNOcJVS
Rai+WImjkx3cMVYbkxjq8Z4UpRQ5ZbIq3+l5vGJdgg6ys6pk6WFCCa/sDqLvpAHOVBTuceMlRhWS
zEEK0R9Nzt3vQbEqjOrwxU6CKJ+6bN7t/zpfWKj50jWr+lPFBKCoohsn06wA+5dSG5qWoT+8XhiA
hjoU1HbPxgHpEe4sSZ2f+B/kIRgWPujOo8dkAvwl/uo7ZbjwZ1JROszXvVzAEafz1wbNcRy4EkHB
l0eixrLEZja7v9dcJvFm/eZUTxKotp/QUSWAOVxHtkjK8neqfxeLO5qzjoAe6FAaGGrurEw6oQbQ
lp52iBoFTq5ipmRaEzN7nLV33bYBmmdtJfpGeQxrWbqNZgYmOj6A1LNxeK4AZ4P4XHP0b/iA3yeJ
lCkRZpKioCHEM+fBkNSfSfkTtjUTdt3mL6fRktm6RdOJexDNx7qkaMVcZ7l+4UjJxjuxlfNTiup2
X0rzYpnn4FJZmlPHFbdPI9fJaKaLHA5j649bVU3iRB25SeSfxZ5cwEo0nQY3T4eS+p905iEvkCFc
G5X13kkm2Gul+9Z72+po0Edo2iWs+g0urD/LbF2RiGFINMpov+8jf1E5WoVxa9YzFnV4bs3Tjwol
HK+q8cxCMpXvdIQD7iciEo32V2BUv/JYoqjBapc775x9FBXRWMzilLgRwwALYDCYwA9TApDZfF5a
ZZ2Q//iXIR7dE3wv2W059X89pBvstkClyPkrDO9x/1G4yrk0Li3/QQQ/94JR5R90vpLq+lrPoF0r
M5nSA1W+B24vCDSEG3r2ilgoiTht1SnKIPFgujL5dp6BoVgSffnY20NIgfJdIPeJhVRQ3NHYNJ0i
Z6CDgIIsGAcgsyEzDjwjjDfZV1BACa2LtF0WbPGTGrzMAdjMSvNTGhU2MfWnWinyIeQ6Gvz/3oI8
PKXeDKKFHy5rMaohgbMRQZhAGhqkbxqX4nCxdmTtn8lCe8ssgeOU0fjKncF4D8llcJoKfqbTfSwa
Rkb3Hq0Vd3tgk5FkhrxcAvCgIhNuzeYTqhCi7+fNDwI6HByC0QBFDLroiLxy0Aj54mHbWgv1NqNj
mFVqUcu9jmrTjt2m0pIV+dby5TWQwtnvbKHEKN06Bzf4LMsy8G7N1IE+ohB7LLPar62I570i271S
VliI+cwMjOGoPzeSqgoPiTcTME5YBqQAL5C3ZJTPcF6wpSCW7Dk21mnwDfqHzjt/gwTsa+8ne4je
87bR29U+5zOrCB8iD7u3yqu2STEeG9TEZ2Llqz4ZVB6KlN/0WucFFoFn7ngtKF9ZIMDDjbUspJu6
0gvx4WaIUlXsiqSLREuduY1WwoOdLYfRaBAL/pS0C2PQ+dVM3wYa5X6IunkNbU9ERGgPqBXwhxud
tgLu0OEVOncuEcGn2jj7P5/GOlUIlDyG6xrGWzcYsdg6o43ncmjkY9eAnbpRhjczZSf+pTqAi9/0
SXZf/TBgntnIIkSakBjolGIZEsU8TCW+lPiR7+L7nKPogI1cl8uPyJGFxKg6JrKFJHtZSf5K8qvG
aYqpZrOvaOrmgruyreTaa7kbcZWEezLhEQ9l2UDo+wJLzHvae4Nly0xdE1k6I06iIRnw2FU2kHGR
PW0KxTjigD889p160WAhbpENbvmyZrRpnM4o55ukTPxFC2Q7QFIOK3iy14ch6q7NtRu/QZd1AugG
gK4PdgxX39GkjeZ9/wGl8doEjSFHbDLopf+ZifMWRRrpdzKxFl5IJUO4wgBgk6JMGKXxOhoDyQzR
617gfikFUyOatQqFlulyAbVSMQA65pjkBrHPAQs+BpHcVvr7py9fmeUnuQAPOW2J9EQTzL/YaN+t
qe/oSnfSIAYAMFbtnD2DwlSYn2G4ilQPgjoCe1GcbRMvoOMP/XFF4mb58/qi0BTmCmQtlhAhU5oF
v2kfuyddwWQv/crUob7aRws2QX9vRFWT5nsCt/2EhUiTcMyXF0z5+dg9l2bw2ai+bfm+rlR6KG3Q
Fhgc0BzGQX1wFIxBZCSiHS4fYx6EAQnm0+id82RgU+D3FvzVBmtwwe3fD5JLNY2ruTPzEwEdfABj
b6EbantMoGX5hczTf9TePrQHLyMdp/umvuRmGQQ1rs7+Mt90/aW1W4L3vQn1CHJHpOMyFYrDa+PY
xwFfcVW0XOogU4ZSGzJ3VcGh3+fJHzgDEQSGXr5j6dJwMJw6mloEicOEJX4oTpHJc31bsuLVoYuR
ePdUXP4p3P7TA82sCH2TW6kamFwEi6VEAWmZsfr/EEWkHdTyTJSunNc6+kXoUKKdOqmhxTXZANs7
Af0F2YGmC7HxJsjG2KXrkGBEw0ATQrensppFV4jvAlXsTcVPX1vB7x5/MndxZNwYG9UJ0aINCqal
kLkEUBKtt52DfM0c0TV9ANahFmwTRUqTVIGbfeUe5EwzxucICzji0vTwMWbvB/qWZtDW9q/RinH5
KFVwBvMuGJYuWj9pFhjOUb4Ud1TcpKWrU6RVs1pkJqzWuJq9IKI0tVUffnuqcKGK/4S1jsuBTVTL
R0sDv6PeuwvG2eyhuwSouqck22YfYqG3mCnM16zGw18601hRcNIuF2Vn2SakzFpUYXh0fjTG5ByM
w7T8WdooOqH44xKdTmogk1FsvZUScKeWsJnz6x8vTN7idkLGCVJgXYG/GI+La6Ed18U3oNHziV6a
xn1a9mECNGm9SUW+xUOMaLu80xAXIw4cSdVEVECxWOqzJHDA24iM8Gmc//67vdlV8frggMVr9y9k
1WmKiQRvvuaD4rPU6EeChXzD/2yk1BZ/9RgORspUQ8Qyc7sDGl3I3C6V18dwtvHdFFCf97N6iSLt
lhRfkfAKaOaoiH7QHwW7lmj0g940dlPsfafkiJVGqpUtWzjxQuBll8HWvZhXI2lqXQmWH8qxNGVG
8H0NAN2z7rL4DRg/7pk4r7W8T3cUIZhCnUKbdsTVD5bADStqI8A6M5d5hr2rziHT+uMt/794HlYa
jkuJmxeTR1PrZqZHl5KeN8fes/EeMlD5jEMKlgUO1pSnr1fOMAEEM5rEPxnqeDWuj5T0rsHOxg4V
1Hjhc7bndcoIdWPvMsRbcAD8Dbo56OAmgewZx5EqL26wOsjejf3YTI3/4RzM26aLR/FePBADRb2O
F7HLX/ra3h4gO+WS0w4ClfF1xkJB9ySk/8b05qfoefmTEiEPWu80dSfi0LcqtVmTbX8Ko6GQrRjY
KDHIEE2U63Za0MuMz4Kig+HQbXYExy3I4miYL1LLYJasqkxsJnf/YCxFTmlxU6+O0iG+D/EkgpPn
ZTlRT/oh9KDuEL8gaAFO28d+nIY2SJmK7w2upi2mK7UqGAbXGBOsX12qKm7IhxcYTxEz9/ukvHKp
+W1cvamupU8N8jaDyIBu08bOTBcydX7Mfa3gEpWQtnLLjHQ9VVzpMBwDv3GEMhXQxJVljbF7EXcW
aPucHyQ64+lM1gKrhK2zFH7HzUVoojRTRXBe0hJlvVsX3LZ0aQPkbLKYkt91X2we0gZ6PEZSdN8V
epthcvmMiZgfWnOSkdegnMPhAWMmiQOGPEKSjMjyO9QwxXy6VDVym1WWs3nGDX4H04NrNodsvIZL
KYfqKh2cKYWU/0HCprzm22B/jGsNkwFHWEPIRMmheY/uiVYaS5p2UGUNlp4oTqILAHpJxuj2Z4EA
9oLM6ldX0zR2J1PMbhx2Np85g4PTLBzNPGBPG+uHbmpN5RgZJDARL3G9H19JtlTC78FnoDAXtxjO
+NetuU147WsYWMzcHvczxzGFd1+4eDy1CD4EGpSwqAhZplhl1LqvGhmbNwdXCWHLtN6FF04ZnLEy
jGAPYInJ3ef4xmnoWkx6cpypMTWWgXz9uZyu4oaRhFNb+PfFVyLA5Qo0KWaa8SN8tQn2mZhZ0eK7
k/LGBZDJ0X1vW7mKJEEplXNnWgDXNaeyl0zAW4ZbUhRdcxcMGKMvOS2QIV4s/jaKa/IfgLLkaMa0
/037rzjAeK88ZOPs0fUU4d2nLGH71eBjovjjRxpAkawnn4jhqFYuleN+mvnDoCLUukr8yB3+wCgg
Q8ambNCXett0F4WGUqr6nexbDIJemyv2WdpOvyOuY5IuE7hORSkeoQljUYZEo6uhVDTNhnbtC6u1
UQobcXu3O+zBxUejT+Wg8cNbGg7Xpbn1BoMvebkVLwIbgjmU30XQGWNqLVfPeLijgSbZcUyqjCqI
HOxmzW8tB6GRwV9nhITlhuOThKGBYq3S2A9ucNIiVoNliGh3v+CTBxvIn7bl/DALvgOkTjF2fO2q
OpyTPfY23QbT4NyA9N7nDyAPoHtS02i3vocPBdsK7DZ8LKFkkwVRwjQ/LD+dhtalyVFv/yQdpj3e
ZrC8Cb4ryvFMWpaMB0XoTMaYyXFCP5pryOuRV12K4bJ0i9nkebru2TOFzQwEvfDmw/Vc1L5BAq0X
wr56Wd6ICJ6pmyw7ZRv56Qq/VbCriKJrBE5Vs2KXOqWmj+YivqQRhakW/ntw7ZzD3myX4bNfjwnI
Z6KPqMarC0J5S06823M6weImVSwCKGcrjMyATxzst+C8ofAPlDaeb/Q4iZDgvNycqRXPws6ITZyJ
Sgizv7pc7nFpvzLgMfh/xBJYtwFSBobu3vAZYff+85/OGDeXA8XwJ43xj9+mjxTSnzDR4oKWVN/j
Y7heRfcztRn+5bi9SVH5r+ek7/Bl9yEDZnE7s7PnPM2jsn+pYveZ2WWwdBSgWLrYB36Dx2TMyVia
WiMCqyq3x6oE/Blb4d86AbjKAGWCO+PiY1D8dgSVlpq2pd0P7xAr17R1uqcZ4ufWIESk5Y3fhwgj
BYuXAzJmvAx+xM1sgnutcpVRTIQrAsABeL1GIjbHtcljK8j7Dx2Z3raJTc1juEOyetCefdYpmY0f
8bXHPQwpKpRow0AlrYhJMsJzqdsZ/4ZeLz+rDR/zA/7iptwe7k0mjzSnRQACiZGtxmvDlVQtQF6I
ACNDwzBg3FKf2vBp2t3b6XC+mIed7FgP55EIvOuC+qrpgqWWQbPOnt2QcnLuxP/RpKJ35Bk6idlT
3A+oLoSl1PVMk8ly8UPt/qI54XbHkQ3cb+vqGbXLy8riR82BbFCZM2QBXatFgSpWO7jnpXYYqw3b
HxLorF4M1Is0Fta2qrbRUTaah6BQU2IXlIBiv2KeJYreLp/D4FDRZnHwnpep/Mn6E+iLUiu0LJoL
0I310f76X2djmq2iitlF1oJahJsAo8GGlcJ31dPy5VrtD0KvYbRqd9hmR+i97pfWaIGYY8dTF7rS
MVllUUG3EE8kGxhQERZkAKPpFtBgxF+bwZnbHFhyUrgoFumnMuP6GOR6XNOhUyxDqR8CW9hwaYZK
gcbvrtwmXJYvlNL2ueM1LXUmWFhwlw9YBXSy29KqPYOdypu0VLKLZeL/85xiBgpBc7nIG0MUUCvc
GP7mvo9vCAjKEE46TJPLlOoElKlemoWghZ+rp10Jmt5zBiamcQhJiBerxeVKu+OQT9aiyC1NhTih
IwDdYKKKo2rtx6FX9So8mT0C2oH/6rd5UY2vwY9mE7BZcXxmZ0JjzqYor0XfQrugA3KE3O0cRWo5
vojp17DlXdgN+qdb4/N2FxdXq6PXvzUw2D21H6lksyM1u3rWk2ObZvkFGUURURrG8gGIk5jOWSMw
OaHLiCFcbRmkfnlXEyKMlfxZMTtzS5B0Rkffx7G/tXMW0DgzYD1BZ40UjZaTJi0jghbGFiNjVddK
wc1AE9dMVzsHQB1oEbjXzND5aPJGdLVI3Mhi3nD7cs6F1ffRwd4zQ8ndEkDDa3XwVMNS/xSRRnXm
I//BIZhXxvZ3uZtaNQsXQI21Hw12MJB0PD4rifFDxXQBlVhTOVxzF3ZCQcEg5EHpVHtRe4llp1Xh
JdkLIksVjgqMvTl0d7/Y2yaTjaSqJPisQeoTaGPom5g4CjcIw28iJjN13hM8UCYcccG4thwBvRy0
6xuN+6jUxwV9ryZglQkzLrgtCl0uX0wMWOrSmFfKkoJ7GLgvMY3Rv6Ylv4H5mb5wAQGQWmO+Wi04
KhlTzahdVsJD0amSzqzsq7l2MM0f6RVNxt4qSLNw51SlsOPf4Ng17l7w/6g9G9kUzx6m17U9kM3h
kmxnzoSVhSq9v1+vnP/Tqke6f8mhq8JVlQzsNk0Ct4AQcWvEGUVLmKo9mYrP0TWmeL9n2QtSEh70
AqGhPe6rD1yfvdLlRMzvqt/Co4pCyKwQn/SGdA72x1uslzLhuuD2te79nk9K1drnh5SwPQ2W0zKM
IBcF89Ba6tLaUC3913dvWoQ85y9vrJdgM4Uuq2ppHYGay0luxeab/8PnMjNclBKC8UPZS7P2Ji8I
arkk7zerG6VzV50VZLwt5MxCB1TAbNqmelpqvG8U9Uw3oU4i1Bqgr5VXZLbpeRvXj0wOthgmgMTs
RpSrUZHs7/9RV6WWjtr660dMfiwLJQweSJP0Kh1wnnzfFqpjSQEv9OTTc6YLqeJGf+hmcemshAmh
IS53RX/Wl1uh4DrPNf2xsr5PzLTiKIC/eO6Bk20JgfVVHZrxUE8cXADXbPzD6sVlWUho8oyrLUZL
FqpR5ktZYZJKJtk4lFEqRdeB2zMvtjCy6in0FJcbvGW+kw3KcFlCLdil42Ue+2uVx3Dm4LVbBBk8
RtehQbNPZFmqwKa2yR5fKWhIZWbP4A5jDstz5fBXYoR2fqafh0m2twn7Crb0kltQIwtINp8eoKBt
zvZR948HfDTMiwwIp1I+s4tNlOA1nLOTa5VyEVBiHqWvoFHIXDz92Humnh7e5VqDOhLxsBk8Bcpl
nLI0lxfJiFQwOP65p6woor53m5EXovmsz4gYrb2T2lQJaPo9wEcB2gyRweXJrujcAr+A+8f7Zawk
+Zd1YhyNrvYhE8WNhRRv5rqBIndp7EqVpGXvZWaV7e99PAwxTV6k46Kiu4H1VUiFzNkT4tGomBo9
tzZkZtC7/1CY7JMdDtvuG+tWyIkW03FaEUgF2Kx5zVgLdS332XcAQ0NLkFWOtfd2ByfpXWXkWlBs
tAo/MqiqJy+BSOIwXGtaX01ZOblQ7r26VlMvoD4HKcSbh42LQOOXIEcBd7kPm3XvW5Aofs7MPaA+
psi2DyUOVjJjQrFkZKdHnPO9HPo++o+jeo9ewalT7FYfLUwH0qmszl9BbwQEb1F3M8ETkzecvmDE
KC7TkCov4DyMIgfcFrRjbjouVSUoy9HQBWyysjhhs9NfqtccfNpfGwlC18x4Il5lZO7mFS3IGLID
mtAVZfJwnP85jg5KVNDH8PVGsmhw2PPwHmoG3GKoVQMRrqwaliAg8yKDbe9icW8ieZoYvJAKInIb
yB/37LSItHblK1zA0ll/8nNBVV4Lwa/5chCzb6x9Q+ibNjaDLNT6DXKl6plwkGnYJiI5BJ9pXlH+
khP177Qs2vRvdhcoDCkYVds4E1GmaGDJQ2MObTrKYSGbDhi47HbbygNTClMvp5U9N45ExBqVSBI7
+yt5e69luxRnGzkeqUP6hOs0B8iOMwCQvSFjWjZTWXkR3e0LKELriX8RcMOU9sxTWYqa5iloJuBo
2E4KoQkQPw4LEDD7pk9QAT4MVbUXCu+YtYr311x2cqSyYisU1lkfzKH487ZGuwBfXyOigOc1a1lo
7MJOwb3p9aYT9mzzhmk8VwQL5eWuISIrK9JQYAveXSRknq61BdNmyLTUNrWQo609dGnw8B5TsgHX
uu9/9Ao9XJmVJ8p65JxTGlA8bvQ/hrViuq81gX/MVfiyLNdRTlDKrNtHQW2O0vikB79HJwFO6KgI
2sWCtL7fIjrZDjrqqOHrwRrvMaiCezgw08guVNyy1OYljgTkkwWypW/DdcUB1FmEGly4bWARIEfm
0+6ELcp4Kpz4dNFeeEwIEFjDw7KF7s0iDijbZ5lG30ZqxXW2uWITPHg6fWa5vsO4i7Khb1twmvvW
gYMwtJI0o/mG6Vn1RM/h2P2v4g34uS0n7GJePzA2fS+eoJSo7a8QOogqiD/cihPZJUdA6uOlbOMV
JlptMjkgd7U7aEopM3FpSqnU95xo+IO2B8Fucqu/MFGXFDaXmPv9ueMeEtMtQ26pNYTNY7qZDOOI
FyR/3XncDvg9O2INIOorek+Rv25Ng/lgwjO7DvbUBxAmK/T9/tv51Bq2qw1jtdF9rp0Lk5iINWVV
6ErHybkgge8/i6tpg6ZS4y7YH4/zbTb6cuPzvxdbmg1AszHLkWjagN8XxqsPCOmZiF9tBP8p1dlh
fG64Q5H/4M6Wiwrk11FXnTRmjfxlQJ8pQ065GiZYjA4OvLLzYqDfVc13HN9pQ9oc5kozbcrA6pPQ
DiYl+SO9hPibBq8WZl5sIvKRgAgumlzfn73Izl0B1YDQUtrOSzmEkBCG+pDe0vf9tL4fL3M159Yl
yY7T4DuQm/s5mGNDqp+uBkP95y3NiX0YVqWcFc7l3kUV7QhQt/D+yGCIpZ7NmJiYVa4NPJxZ9zGN
0402ZuTbAjkA5wy4riNsoBjW+3sjBiXpx9Qbn7zOlm+vs9GkfRNitQoodjkiJddyBhCPGLCrCrF2
qhaTp1Kcj3psomi/17SBJERVZSPOUY7bJqWFa7OyEPYLDYMkYTh7AaMBMHxacepV6xUmRsBIULtF
PVBCj4ithL/z3y8XyPiyFhNzAGoIkX4JYnQQjjplbHAduzItWX/QNMNBoMwPg0gHn63lBfugV20H
4MCy+mJscO2x1c2CUquUvbyBgcI8T21edue1TqoC24PwUCfJZc5OoP4YyPEp0DioQdHj+A4x6HRP
WfQvbxdXM+mUFUj/o0i+7Dt/Hzb1qNcva9ZisXusLsf9nwVwErBvCS3xBfw2VsvjmCoxV5fAN5yV
zMdb/I4HL/s+CcYvpq0ny9uRHP2lYTXUyJ6os5hS3D98yQqSEGWz+vpCpARLXfEI01YWgciaydK9
d+236ejda0Y8h0Vxg5Gi6H8JspiYCkNg8NfmIdA4VS+VibYggyxf14CmY9hUY4o2hC0b2mvDAlTr
CYxP+y/l0mrA3NBOjY2kNLsOdTnhc7EjmdNy73wMnXvPtDbbDY+y2NYhCwhkvqzTV01pC01OXf0p
Af5fwr5NfOCIM1Y/HNhqw4aDHqLyeJ17nL1Ilkv60k5LLh6PonyiaSsh9XSTqdnGOnoLd3ddFKSR
zY0/Vo9Rx+ILDiYISx2JsGPXNGcDOUUDqCu+wwOuI7wFhedSIPp6/tBNjeyr95OGDGbC2h5GP917
Sglspgz+QvGDdNI1dWplzn3ryXPZpP3MR6PMtCGCyPJwn34FzDlJmlf/T3t5OJBwgO/4joCwNpN3
K4D5CkSOhthvG+NaqHoGqYKQD7V14+WPSi+KutPMA8l9+Hz+UM12CLAgU0sAFIWkSEckWnkBcWRb
XZybB5i6z3uk1T4OgosDSNNTKLx3DqWv+jey8lECxM40NJxZcAFyV/VQ0At2tOeHzry8Ky7XyNXe
oclGig3SJSfdplB59XiUOjSGlNU5sN33mOqHpROSv+aaML75blk8KeGIkfHzK9Pw0MyHCNEJow2k
R2K8Q0QfiDM1iI/Brh3YQgioRVEE24uVXdSIukq410tIf0PN6SNdbq6Kg1eW9D66zqiwwY3I2Mrv
OOMswIEencyqSSM5GHaHO0vQBGQbukSd9XhH391ft0Z+4/iqd+XeD6CYeA9UYU/Nw8HoOkSFhE7y
HQy5uwZBVj23jmya+6vGVZg2r/OPWC+ytswjQkH/5b+BsnpkYIiZZMcILaQhIdpUB9W4JGXMXEPZ
tMQyNavf+fevqevr5pYiU9Tk2rm77Ft3dk3sPztXgrx440K+6QZ90QOocSI/M3HNI2Ynjh2wdQCw
uvBU64FDiQea7cfCN3W/6C7zQDEbsOowQV4yC5wgM+UWj/GT2we1qjm0pPdu+3Kr616CKjCzDAAl
Cy2ea1m9vnFrW2yk1nqPTpK2IITz9nZvCg8/B907jlNMnsQgGHDJGvnTo9c/IETY6lL2fQ+tGjRy
itH4a92+EPc1TlCRQKMiBlP0dLiv525NVQYmxvWiNnqy/RE7kvv2Jqnnz6iKqWF93T8pfIMN4eRN
Ll2z0n1zF3Z9tMWxiF148rMhF1ZyqYkMtYEv6RGHhEMWqE4tnuzqwlr8DWsES6d7bLOl3MjvKOgQ
jpm3KwaiGgEbE4DWD6pWhu/P/VqijyiimMYecn0Qn9ymKvMy5o6eztYGnEMhbVKvYLiJDRb72ra5
jOD0oc4MvYvY+dhoS0bYDiVt+S7oUFGX+h2PD39XmmO2fAIbL1mWKL/72CYv2DfZuDL5e0rDPCBi
zghagRx5Jb4DpR0y82iCdH4kZeEqE3udsTHkNBnRJIYGIT3JOh5nx+Aco1LzzUlWBZdOGnw6dCHz
UTyWp7RrScSRF7caJSjAcXRArIIFUCkXG7/oQ6+VUTmQQqonuxNe93EtOy7h7W55L4Rl0BwbbfJ2
ufTc2tgdh/6IIQD9e54feQRJ6jqecvt+BIOE5VzTnCVtT4zuJqEhTeo0QKcQG3I8ROWt+YKlZO66
cr9Mba57+oiZ5fiG0CWhxQkvImCaWqUShhGCtqNsgo026x1C9hf1jUO7z8oKQFPwxNfphGA31+/J
rBJBxnX8LuFAL7TrCGZ35aHMUmF3CgUd/lDcCrVU2/KxZ2XptuVMt/IDsxHiiLPYFp047z42dNhc
83H3W9+nnXvRuUbRFnaovZCtuZf7KjWf2OqccAtPgkJzLMP734/F4q8POaVT1JHocLeMUY+Urxhk
XSygCH1duVEBbA4fJMhmBqBnzppr9QIQ3HqCCAfRtslsTGncCtXr1LnOx9lWgwjhCHjYK0Jeoe88
74RYWet/tG8QED4hsE7c1D8eT6LB/huMNYRfBH0H0MflO/oMr4xJIk/b1+vATZRzWXNm0fUpuFzm
ZX0O2SanLYdMwivxEbTgx92KJuNsERyUlKEmBKacoAw3ic71hnNJQ2j4j8dSAVQy49G4sDA1Weda
S7kia4QsMJYPceZdm06AWSzRECTUMEhEahl8cr/MGdOhyXcZ70jN+x8JYAFxwkEhfYPzt+9yAuNX
9oW3Qa4GUprICyPZzGmNJDLBVuHDWYRS8oSqH3hYo8Xx8QExibUOKLMnWTCetoWfJM41aScBESMr
mAD582af4KZYQIwyZAUi65G3kTdHsJLblGgJc/pdZxMFwA72bXxHGnmxpCmnpNYu+1QGz0duw/8M
m3zF1FTvN4M9/zI4JVGA5zXS05vcoz0BkxYMsKxwAkB4NY6PAPM9+Uc4HCfFt9jVcNAvySKCOD6T
4MM4aO58b7SW67ClKgskHCE3XLpc/7QGX83spWpm3eY8eyCCnsgJu2lLFT1Ehk38H/NmZ3g1Rt8Y
H3PsIBm96sic5C503Y7votIYG64qh+w2JdRudjrfPcaXt7MBXY7hI6Rjw3K250pXxs/1qHgXHYUZ
xVpI59/cM+8rNdZnZQiStnPCnEShJPF/BErGq0GbDi5aB7MzHySCdICenKNXIXW7H23QqTZYJRqA
tUUON77wceJASME8tSo6ao9JhnXDp11aUzpymz4iFQQ192LPPPXD6uy3sKpOrvc2/RTqLqs92VqN
lDrknInn5fYXicKYxZqlRYa2lJrIQm60BZ0TEbhqwANvM5LK4+SaY2JYimgoJ1gc8492aX5vY4JF
6XdezNQSdTyjiN1lEq3uQxW+RrhsdBhNlbuj62R7uFBlIkeJsKhBH9KTap1pZBQQ32k8qCsWzSzz
pGfQZOTjc9Hrm+L3zelJKPnU5QY300C3QKE0R6RsYeqagYa5pxoOZxR4VvT63autLf8Yn2nW5Qpm
9XSI0EAPql1PWq8dCCVU5vPe5WEa9yiM4lmZ+JWUTwyGQZnO+PeyuvfJynnDY8uNJpDvZgxOcwDB
bPY9k+lGB5Jx2IeC4SjGWdy4rjxvgUSTzGSyoXvQ2ClU46gH4YRyxQrwpQeRdh3Xyp9wTDLW3V0v
KpiOam+vxNvTJvIQSu+Cv6WEuuUGK+l/8KPxwTrOTr+66LkYX+oYVxU7UdLuQWs34QPh7AMb2tGx
F2Vl1Es0DZZeWtWPfLencIVpRCtu9MUI5pUlGHR4Qv8f2Flht4bvjnL/69kIEaUB1CY4VBna9rM5
qNqYtj2ydXzamP1YPsZ7tKQxUjmQ0Qn/0R0zuiGU+JKG/0mq+zZ5X6JyN2Pdq8qs8JhgptJRs4nD
6kj4eEbS3AKlrRI5hpZJdG+B2+umg/1z5b48rcHVN5iUwEpJuqNIwkKGAXZfYiYNyipwnX++dvI9
qhbn+iC6It3XDU2rXkJc2M7T3QVjg+aVtQe7DBdkbJPY5PlK6zuXDC4QYoTwAVaAiCd7moX70MV9
Cp90gmEfjU1OYb5CxYx0ERJHFmUDTN+U0g0+qPZAUWJGGUHGvtxCfAIqSQembgLq0YTnvpENfAYe
Y4BDxjUEyuzwXo5tEzF60Ea1Xb8/bDW298dRJe7NNYXPbf/a+L3dlXZU7hVyWQUSgSHk69pHwLqO
7XHMuPyUkkvYgAeZ5fLVElP6+QEBQG8dw0MFZKrUSCBNLMkOM45s6iUFRAWRPGZIvF4w+ZGr2YOR
XLNDbbBY1SuARykc92i0Xq8j6EPcHOr6qC48BnQlQ7b7nGTWatgyAwzqr/pW2fWrRvia3XEOjXgH
qP0Nv7UNPBLVqFoHTiFMdVjHLZIHFzaj3AjFDSJsdLFel5cw7hkSFwDXTSv0ueAvB536pJvSYFoA
JhNOxKKDFntR7z5EgfFv9t5zozMshVEIYO1WwFdG4CpuwEB9ed2XlFd5gHO5HybOqI5k7PbSawKE
GwDVz5Thg7EASKHEvrZmjxz8DhEsriurbPXZ+9HCNITWcv+LiivkRatJYNSC06iN9LVWfGmr9DC2
dwnLsYFw50YvIFaRrxPIVi5aVaNMttMMTjzjcTGrU4VlOI9m33oaJGMFDQVMFwWVVfI87PTwVkMp
JHKNZGUdqskGn54rRPzsczaumoudz/oOipDKKqCvPvHrd9FXrKDb4mr7u+nrI1rtI8D4MnqavBUz
h84OibtOWqXO90BQOKcCK/qkOxvsLAsUH4Ol97PoEJihSAGUf3VeLUyI4t3hsclg8mOfBlgwtd3K
h6+I9xnn2NFhMTXE6ZOzI62Cz9QvTw4WXtHXrB71vcKu02QymfClth42JgVNRTbREecniHBNm3hE
Iv4Gku+78JRRiMuNNJVCbuIAYG0lMwDDzOsla6s2dqTudchSdE8whRjkMLZn7ubhGWuTdJydD2Je
rWyTNrfexnWoI35A+/f+kPWXry5N/LqdHByF/xqxaFnZYHvCPa2jVrRU/GrwDH0vKvlsHzlyBOHW
/0DhsLVz9YalS/LhW9rPyBQSHRjMOn5FGRx0mgn/txzMnzjsbbdCsEyQDQrnlk8Y2z5DQVgq+HXB
bXTW1/ZM1+IkjsJ/prRUpJ3oQc54fWtiZ2Np0MJEj8Y+GmRbq8d/IUN2k3CDPmpT8fg/6EVkS9Bs
9NJ5pxH6NyYjqtsGz3l13a4ptWIk2PTiU3QP9l5mIYBJMyXCKjkZV7l36bXP4N+wGC7jeMZ39Rzr
bUuxU8bZUVidXwuRHx9heded/lHwDk4vx8ZgTNGu2tEBx+/WG0qKMDnfk+2wcsD1HIztIqQESk8N
Jcg5Ajmby3mGwLjiPpQvGES04CBnDe/U1VdGBOPLIeuxfvNBmcDiZz9jytuXRW+ixBJMTvvDbe4f
Fi8aSw3gnr1gNyX4yTSDOJ78cm/Oc4EAy7IjK6yEL7ivRygovCVdC5icZCi8WZivNkC9VXi21j+z
FNsNsUEDgAS0y0xK87feL8JSHv/ResDq922cGTlKlUdzF5mSRCS3bdam0nLY9VK+pGfHhtGTofq4
y9Di2gNkPyzPtKACRyb5ErGkCUAA3W/vMlIJCDdxaq6HSYKYC0QTnMx0HSJjrhIkwHjvkeroe7Ik
BeGDTUb+YFqxNYkQDmGrRpJj/SJclhRttUz29eJlH9eLW/bSTRKDjE/TO+TD3gkDM5vie2Mpapnz
UH0Hi7Put74qWyiN8gF2aqPDSfA3eu665juJEmPp/0JrQkXtV/2i1dj02vrkhyNI8u6y82kKBMoO
X6NKM2Ky6zwVquOmfr0LyfKdPz/Y12t6JeDvquY6Xram0wQSi1BcpsBzo2tP2ahMUpf7msOxsD8s
XTxnFTBdyXHunQyjf9Gz+d5n03Kc+D/I9f2neRjVmwuKkgHIL200xjaL67z5VCmGK0Bv/xTlOC3Q
EaTIhOAsBn6NH1H1ZS2QJ/V8kI8eEfQpwKAHUhLfYPJMIMiW47YzCrg8aFF1lX1jU01d2cvl1yWe
GJZriVFfbNy1rF0OFaRS4kBZ6VVkfimWLd26J5gBnjnXCK/NqzdKJjkqjqSrrFE/TvvlQghiKv+D
/EIFFaphQkXe4+CJCt6xl1cbhETT0DU0fqQMxQ3RHyLpfu9S2FEhpqzXJm09vZZJS7wGTnc3kzLn
AkEU/XbkiuguUgAW+tmqP4AOR6pUbm+0Ce0roZYxQHp5Qlx4IMx6HMi2rZsUhB4ZtZzbAY47pZuN
Ti/3bBGGD7Xy2AFLTET6mwYtenn7dUUJRr5WnqO4TG3FOxgUrz0+QksUNAlHrVQIKEPXxOtFlo6u
DsKqD3Zas9n83HqNUwWaN7MlA0CzcipY4bSHvWOJ5sIgRyfc8+l3Tvc41ou5SIA5MWs1AZKWQ0Wg
bsNhg0hqrydktWDmPzKW0ixJ7DMJa3V2x9awzYvS4NaFrbkSz7YGDpXO82+a1iWrripg59ut3Yeo
qBcKySERuYBMQf3r5d3rc0nDxrEoehr0GwR7+TRqMdEhFdEoCCO+FSy7Glv4kEoW3mLHIrPS4N0f
W587CUxy2EIN9fEFAZr8yMPXXUy1L05FSC1dEKUTWJDIe5JjWwp69eKfduQ1TvU3qu6qL9CCCl2v
SXa25NgS/fVk2UEuUosvUPxoN6Is8pynblKlbEiWJ2C2JqMfvhJE6QyovKUq7vWMT9QCgBCiyPzc
+qcdRjg5LivOstz9aOeWpmm/HI5hJca9Dv0kOgn0lpb+DjG4shsvs/fcEs3FCbuBdhE9vGtLTV1W
N8qvgdGq5JfvVKGwHArtlv8m3P48W7VJHjg2tRVpJfZ0Flk6BxqcRu+hNA4yFm4p6khJeY3TRqkl
2/M++Kd/xiAy1KMtHf7Uvk056Rc2iZLQYxXHm8PtZGQr+/o6EBFhXXFiXecDWBCCBLS+BjaSnXSU
KaxYjZ9Ng2LzqygFFqGq6Tfs//3tbqLtBNM2Jw4XLYliF/NbWRAqPbZPpqj2YROwSOhHTfpkraQO
PB4FnbhgHCBYQ8oWn6JXCD8EBMXn/7U4KIzJ1bul+ZPUCe1IRNhhYKtqAseYXvmoM0XTQqwVFtWo
eHGzhvrm5oKczNKEacryT4QMzDd+pkuwJhVcaI0zA5ZrUMg8cbpmzM6z0S8oTDc/J2ix8ZG4618I
BUpO22//GNRo+8/klQxFEBngLmi0WMxYxDSskSaJ6wPGodWaIEvzURgLY8KG1p+sNf+WOjN3D9Ls
EP8xK6l5h0J1+/eXLWcJMjvynxoU6FRSIWOJJ65qgcZe3hWzKFmPwjuTISP30FsasQUwkUcMuQiS
7wDJRbaZ9E5/O/rg1+IUX8eLsoJjOu7i4oO9N/hxz/D2eCIVxdMACUcXiEY0zEwORDVjPVieC1bN
wk88uILB0d+bPK2//6hSk1xpAg3xxSquUFV+MnaJLzKYt14MmHdTlDjQ8cUCNDfjsMX6vKwFUlh0
kfdC/1TjO6Vc+Zh8UBO/7YdU+kx899OeYsUOifXskZfE3RpPHzM8chZc/zuq1/oB5L8PLFgLs9lM
X/RYdcNTYPrEFFo6fNHTW0umSEjtjOv2LVeMMGRbErN/xG16AsEmNkkXN0CowAzCRN01e079m5NY
6XAl/AWMrQ6WTvaw1oIG45I85HBMW1Vgw6Hd86pkBscfAAIIoQN0ta1OfZg/+qd548fXpdvlIgKF
mVJZOG4PlyWoue33b2yzUNR+NdNzTZdAXgx2jdWVFnVtnczJDacTnTjgYaH5zmSo9mduQ7y51Bqy
MBzeCnAtPYNMyK3mHDK9Owaw7MK/ekQSdkWEeigSSr4Tbfi48s8kxLYvQ/rZz9vxViIdhO/mDc70
9+m7nVits0Wwc4UOFrFeaz73FSnEdQzD5ItaOq1BwR9NCG+1ZKCIKvsvIyP3laAuePujimT2x08O
4J7LNQDQkI4Hiq+FpQU/WP62k4VTxyr1shGtkbtSXHPjaWVkbP+rRiU2NpqlNd7lkSPOUDFgcQS9
/H4a9lohomsF04CqVnJfeoMpN9ek4BFkUGdtIOkJIdm/PvpspTvGrlDujvcadBOwcR6yZGifD3TL
7oDDSnlrVe2y+LtssIRbOG5hSNLWu/EoMUfXTPa5Zg3JMPnxs2pFHYpSw2XnfPB27yu4K6kXBVm3
y/bAmWtPJKduUMQ8BVQeeXu8ZE8msGcD7XFFvGI1l4fPJP4BjO5zqolA8XKJB5OeG+QHba9HRDo4
D2qN5epvHIaHAMDJS5RbIUgYFKxi0h7jDt+fR9vSiMH5r1jypPbnMPd6gGwTgn3lwM8/uSz63l0s
gFOGWGdx6o6H4j1EzOcMxpAxw5GeH+bxTjdHCjolcTuaOtUMacYOu08vq+74UxJX3Q3O9O8+6N9v
Lf2wqYcU3F2AAyzfkAn4MXgdMwvL5qd5al1V2knvQX+1yEvjl4tAg2dlc2N3sWxUTYQoT46OcB22
+4njqbXWMGoRqsb2clom3mXgXqgEsAsVQylTQibYGK43pZN4KQ03bsPawRZTmZa6+PUwSC1oTMZN
fYl/SAnZGFrcZ17BTKEzIYUDcfDl8cvA2I+6INZYEtXOCA/TIXTmWoyzmjOYd6aN5/mM+ON5rXQS
bY+54KnokBti4GUUPDMiqgmm0t7vpuUuzfysgxsSzKu0czfM2zDJxi58L6hexyTPE+D+OE88dcn7
oFxhoY/1bSrhSlbUB6pFV8+irb4MFwl+SZ95XlQiU6E18f7ymPX4KZqPVJupOVfZ6Sx6tRrCr0Qz
G5ni2tXw5JViKS0Fi7kstf6eveerFXRUtbn60yg5FZpCWNteWQe/dRI3O3ZhXESV4y2uJqOmv+xW
5rFtBicqFTVw7aM37gSifP9b0nQWJw9NVkPJm+wIUEXNTS2hnpsM0Trj3RsIIf+hpnGGsZ5/ltgq
3EBLN14SCOTbEtzu49MEuW3QrKA3i1C/pgAfOe+TSRfLHj5kIpW2E09wkLjbqGXURb9XGDyAnE33
+kTUuPeVVRZeghkZ0ULlxbA8o5DRg5apoKFjzRsPKhewYUxwMoFtfvjNUl2lX669xjo5zgqU0Zy0
Q9LzOMVE/70QQY+DEuzpalZcxwgajOIsa5I4i/G03x4jEbJzgaprPCuFLgovzBj/+cXyDR2wP5x9
MgKcPmoyfX5PMm7MqNx8sI4Euk0u7rohhmxgeDUjsvn/NhZ+3d6vuwyHEgg2U7m4HoPYacgh8d2T
zL4MrI2zyjxI9vm7H5C7Gy+zNNosgjhphcv8OO62+hIepBZgH+mdqFtspU5dX22wdFiO3P5c/tr4
PvLCUMv7sSgZqqHYOpNOHM/0qfGwKC5ZlhA5vF5djXIyPSNNMSx57n0dJ9EvWtITH+Y/WmPdf1Wq
4xlvNMaj28AlZU6okxILRO9FWym7dnCSrPV3psZ47AJKSNKwtCrVTaWjo9RY8zNBzEdFDHmi3+gz
RRMqc+AJLCfPt2hE3uBFUeM0Md9j2Hv8x/Xsf3AA4udG8vEF7xg85GRdKKupWT9JYEL+k2jmzThr
NjTvy7piIlx+aVOShkNSmnfZBSZhpe6naa58JgxH8W8pd+eF05Mjy4IR+y68dHRi5gcgs1pbPFUA
Mf5W1DodklskeWvnkGNrA3BGis1iuAI/rrKpnLUgrt+aqHG6/8B42PKqiU+st0S9UFinkwQZMDlh
19ffkpcS64tB2faKjxfvAV+/GoVZb8o1hlBIp0EZLZcXjuC492WSTnZu8ibBsSR4K4doYR0tKHu9
26prxj9hwQXyIq2S+tRcZktDFNyPcCnLnDTyKbF3gjNbL21ak8YXrgXiuZuXGTrS2+TwOC3iMuaw
vlwNlGBkuKOo0+MWwFESbQBFc8Ybp8fVNza6/NLNzmazKxXsYP5TnSI3yYNWWtjvqd4evkyEloQy
Fl17wADz8ulgKptN0cq90Ihe5Md0mNgwj/rQR3J8PVPyK+08at5x8w5bN8dBC8fGkXs/gWJXUXN8
FBk9/4J2NTnEI87Z9R/GITyIMYvKDmcZdlZWeGUTWkagtOGghz3w9WlPM6ZyL+ghv1cKhJOhVmj4
XayoNOaIxCWThwQ6y3sStJVRMHtFvBdi6ndwRSH7fTv4APW8pdhvAgi0RiEtKqJZfXKWHzzQLe0N
YrZzLudJ6CtSMbAGQCO3KPQt9RgQU9tEMsMCJ3tRgjynQUch9vzhB3nfZh3x86F2oKJrJbLvHQfr
98/4LOdQus/x5HHs4ibnuExCtm7TVMSE1eytOeGS/YK5NGeJap3o2b37sGuK6we82LhHhk0p2g2Y
q6kJV+w2ftD8k3BnTuxUNYsCMtLEDEg1Ex78GdtmOyLTj+PKTjmOTtDgFLoJsPJqoCo8jBce7lOT
8LaPDsiOb52XqVnr0EgPdoBK4LpHu9H/4unoQzLt4uV4wNAWc3oOE+Vq0v+cLkyPxZzzJYBgxi85
oKJTpWCcmjKm+k38BvGJrJNn1ouDukCrq5KsFs9mqWrPhj1lroZ78fRCacxSOB9vOo7R/WVj/iyw
agYNuTTeCq1OKP1X/64BktK0bZS6Xkal26BU+n+kT33FIVOzP6g3NwX1nMvngr5cvuMRHLtFIi5Z
0C5n4YG6MT8uoNppCoJlO6l4ps5tfShdOGdGcwavOL3M/yJZVW+OoLEzXPFO1kMHlh64MB0iSK28
l9k979AcAZivN8kkW4bzagJplpAqnoON4bca695ckvjm3BV615OYO4xn6w4ijoPTFelahKYPHuos
k2qUcSSSaYOWgJWLEGC/d9SP0mYXiN/P/3eWS+urh7XmigZ5Ik8K1iCpPvGMLtyYMLdlJOgTsl1Z
wDLhrVvTL1HllNqgh0AdqCj4qRDXisBw+MelxMe+49g7AEWEWLujwlhvyodUjXakgZ/zPg+h/eB2
unf8zyLrq021BWZAQlviZoqfFrVWSGsoKPEAKGDeg6S/izBDVZ5onT3Q6A5trSZ4fUPUKSZQMi3R
h3K0XnBYOIbRekrIhWVv6MbZw9MJrFhGkXwmmBIlQXCy47NgSQmrLXXilthmHvi+8rQ8lFED3f2k
Tm7q1gXsq4YU6SbR4b01gHrSNHOWmmMKJK4Xtytxsj3rCKp9G/kyCgxujNtw0ORNyxknRn0AVv37
wyVuaFN9bfdG+rPRhpkBaD4fc/w/S4jdw49wGWcSSLTOaTWpUbH6GnTmJEoIy71buEXE0ACcZDQj
NNa7GpDqoXqJMLIDc7UCerf9K083sHb/glYkhSvwm4JKf8CqNsUSKp94UAhj6uGrleamjt0i81jK
jlVQI1NBqMYlM475jAdp65YBnNxPrnDCIYEG1a2Lwb63GvAlpL46mqNzdQeVrlpoWURj8v8zFqSJ
6A2OiPDSYksnMAtQIpO9/Ha3EGxxb/9DcRInoL9W1O/EgpxP4zXlesL+2lmWS60VcHIDdQvNqoyx
SDmKJgq2BnI3PPzR/Ygbm7bLC8AlbI8654MF8+aDFYAfMHjWnOJaFzzDs4aYKms4kujx6KNUe+IJ
oF8076EdproxcX3qxOEkB8OV/qw1qyO8gX0uxFDhtJNsiesoCTVotgphLQ3pHVA8Ij+fnwcJb4BW
GS+y+S4ZzTyCNp++dA2dvVfe7yhfHxkO/fWw6TjwYna8n1uwaaKJwvwr6eaRlm6kIb/y4YP1Fzn5
YFFPNm74mr1uYk0ktk/TpvbrDtgDz1fQivElTuannDYlXeU91kz7wYlkIV9ZHSdIEFGHz1ahT0ZH
59MTbE8dpmVoepiRQDbtXX4+uJmoDWU4fhATAPFnvCSdSnBQcSJv3qd0WyJmE75fuWKhisgUXl1W
BH63SnAA99Od+ryhTy+go9oYomE8rq+KidJUFEbeIX7DRwH2DD/fYcjVxTn5pKxqLzHCEI3dFffW
1boa4rqB8voHC658MLVmsqZDfnKHIiDr66am5cW+EPVfbXZySdLrNFmhTQKlpT58my1gpMCZoFjS
T5N7SCiv0F/BJsDMrNlUriM+pq/zDLvWIynbgnjwyYdJfPyV7rP3Y67PkGwXaR/0jJh8QSTUEpAs
zgoeRRi9+cxgy9X9XFSVU2CS1RhDxH62dvBvvlfgpACwk6wX7GTKcFpNM5g7ec+9DqmZhRcBC2tj
xy/BJ0nm37SA66z8MGfljg7JN/EpFzV6qDYws9HPgcOD/Sit8jQtVQSV1LNxQXy/o7OP2tosoROs
DVQgcyx56SQeogYaLdaUYAySiCpn6xj8VQtRt5jQE1AZO9Ve+WruvZ0fBgPwhY5FH6SaKCCvaCP5
VP7eAX6bpn804fEX5dTOdyIHd3p83an3HIhcOuFBiA88mfCe5hiStW1VOexk0pS6iFCfjcqUVBov
HZ9sjC4VVdI8lBHKjCDWn6mk8kyqv2ysVtQKi5BXHYXUkVb1GfEdlDufQn7++iFB+d8MlTp5haph
PXK2YjVxxmFSmUGiIA8AZD1VgWTi4Lu4zGd/lzS6+mlfm5lPuqRayUTK1vmHLa4M14ldIHijtpeG
MI8qwIFA0LhHEs8vT7N5thaX9bIPqomccwpya5dbag7l0dxPIfnkjcOGf1mtRoVl/MkpxMKVvauG
Pqq2LSvFgh0jvea8ZYinG0NBX7rzqetd4vGhKj0YIBuEk2DylBV8+6RGxJUUVltSnwBLrPkCh0QM
joMBquvKG5gqClRHRYkT0Qvti+p6PtROE0iiEigiy3B+deNgsTgYWdsAfqSL8JGLa4Lb56YZKnyv
frlngll4hnO8s8cmM/hI+YJmZrEmxq8taxKItIQUtdscleWvZ5Tlf7CNQJMj0xqOZfQYnzZTwMwJ
mEyhww1D9Rh25XkN7X7QYiZhl+sBvSJs56q1VlrvHpJzW2WpyITBnO2QGpB/9OX6OvGX64XcYd7Q
ed6uHOsc2HqCrKRjnGtP5I6SgFJkak+SvmeYOFRjji/lo4yuiRsw+AmLUcfxNtTNAKIsTWC9S2R9
wyA3HBIDzZNQlLLpknuiE6dDiGytsG9wwyOP+gplq9ru0zBquT3ErbzvNoe7CeTdP2f7O21IeV4K
AybO+bapA0c8NIBmCg0Pu2cWVOeWNl+rMPaeIiZq9fQItGEa1CXhpGUz1Il/3XRVpEaSVMpPFkBW
xk+Obzxu8NAK5mNUK8+ZgC7ExeqHtK/XORi8jdYmh9nUXn+V1H47V9IYklxpsmerAAyCmHui6qmQ
37CMnhUhD1u8hNAWvbUMgeUTfLbOuBFQCwl+vTlXPuygWIc4vJCrVZFCQo++V2I5tkRVzGzhkGIT
flWDfwJu/VQIikV87qH1gfbG5TaLA8MAsp6RijYGYIlECioqgyxXZfLa7wTpTl3C0U/yDUj6jvAl
cy0AjxkCYnKJ7XLW6QAseVNQenP1xgOoooS0GmdICB/+c7oKxIJHYPjmPboKgY/kvjR1TrF2oWb1
HSAtcxRl3/gGKUuMSad1HbLN9DGFJCHiF6NBCfKpzlpvJvcH71CQhaK5WfuuIXWlK6Ni+WnWR0bN
ZZYud3UIPhK2ztP48KRjCk9zDvhkSzKMIgA9TiQeUzyd4AjKvuCU3mQeuV5584Oi7hkZbiGs0wGt
uCVXm96nzgCiOdW5p4BTheoLnRWdpgrWWdQ7GKjpRFzA2ByHQ6kOdnusnZkBu8TgZI63tFHmKiVI
y6Mtn9HyYQy/RAtTXfZ9XWJdMc6c6ykWT/YtQ8wlue0YW/busHnlfU8SA0d9lHtvEmwiLUCKII66
7KAgxR4Lw4qfFiXmv8HDjewRG6YDt8OMg07VvLUEiJT1jEFBXqf0ddPBIPyWfUsJ2V07wMvNbBto
8Cm/8O/hWBGYWLecbOG4/ZP1qj/pPiAUSqtQL8Bwb9ZpsQxegeW2qILn7UmHUFOSq8tbcEEF+p+U
i7y5Mur4g0pULE9BW+MNDtrfVkSkr0FJNudsYkbRwxCZiQVwnJK+IGeZpa4jFEABccq/KLqmHsC6
t9BkhAnQR+nzVV5rNIqk3nLBYMzIz2s43igvm0POpgwNMN/rbJl9mQteKaFKF22ZC2ShCZqDYP4i
4sRxTeg1xbgk1ihLGvgaIVKmOKboB45wjNhnQWe5Hc3rmOHxUSF52LOpZrV2sOIzbjzUJozVCCkm
UQN/UvzDkthWPmwvmON/aRBHCGctcxY1xiuRhVlzB3AA/rllbpQr4vxSqe4E+Kpx9HYHMq+cWu1i
CttOcz8b6TR3Wij284jUmj26+K+hbUrpYNYsR481AT7DD+I2Z6QBa6HOxgZnpNSlenpM9MgcvEs2
lkQtbJFKUEwnfAn6ONZBEkk6zHwY7FvegQYhixnknSP2u58CrOeE1v4TPR3/D8ciOg98uSAtthTI
IPa0lUQie0ZxoplDuZ+gDA15e6ENmBRQdI1pvnO6ZDrdofL3q6jpbHA4iybV8DPEKXYtP53cXQDh
f0XyHf4nHAxAD4NvYXhZCYbENXuSjlyMQWzaPxFFeJhviyPYGQTCd8PYrIefn3+CXSVJ86AE9nBU
E9Mx4t4J/A6KSdI1DQPDXlhMD1aNyIB8nmmUy3214QcNtxGCjVaFTTg8TldH0tBcC1n4IvP0GJf7
QYkDqjPaH1VItLvzS0d9Bj1eZ44GnJLEECnOiQ2j/HRy1dgahY/6fB+KZ8er3C8hwnawO42/MH9r
Un/dO0ihYFy1q2yUmLr92KAG+sPX9KDnfO83QQqnGT+z10Bdy2H9JtTIy2kogwYPORj85ZT1opxV
5u6EFYl0S0De4gYfMUbSKRschQnK3AGkytBn4JeTo6e5M2059jm+E2r2GsezaJAX+MKJBu1BKQjw
x+d815DN5YNTRZ58gv7JOouGK64u1qvdS3oXnIB/Xm2KKTnUvxLVA0ZbN4RM8ZFIW9EdW5BT8DCC
Wd0YtEGVIW0I6ZGWSYOsEL+3ozFLjGYrS7I4ONGddHxe03JPgyIlgj1gbbvOBXyiA1CgTPkbtPwM
E2g+r6w844GJa4T7Dim38gfR/UPfKZ7QolxMHDyMvBwK4fabjvVoz3olQO6uqOeiqyfoWMCZJ64G
f+/mhGfX/0g+agr8hLJYO+qFULmYw7Pq3nDjeyK5TbGTpiMyQYZTj4oOtzhtUik+939ideD/YJoi
epnBbmIN6ZYZwRgPKHVsOatVeSHjNNGzegdRjt9AKwRBWRvL+xXxrBrLM3T42kfkiQcpbbLrOVte
VW1S1+4UoeJEgUMEmzNLeZv5E9qGvxtanmSRhBYsMQT957XbXyomefhH74eAzRRlXghgYUMWkp5c
bgCELBfaDzaTMQ5ZWejDPYCfyI9u7tU5vvN6xNwj7PGmkYjeuR769ZPtXenKz9AqIdK5fpQ7ws2p
cYib9K8O7cDBDX9YIA1Cjxo0PeRJjKxGCAtZljNBSi6ia8yl4wDSN7XtG65D6BzJhN1/Gk+gRB5W
GewGdT4vDDKmStFkNUJ/r8VcVUDZ6VBHNaoAcDQyxQ5hix4jyIofGE4CIC3Sau5Vn3d4fZakHw2s
OmTgqOvTuoJN6tMcI0bUvbk9EWGS0aFy0OyBIu0ENDGGhzqX9ceu3vq+nFMLe/QMzmBmly0oUKWg
xWQSveUAtxGD/g+hY2TLRZECOTYd7ZbzzT52CmSR6sbv00uliR2hFFlrOfdacbrdmtqcZ7HIzhj4
nVxusG/Ahy/LBzFLei6W/oQOy2qFMfWQVCSZwQ36bV6wNq2mquc9Q+lxXdVsn9r/ErlU1voFN6yp
O8O5wjkJ26FZVHrOs4GICVFcbk0saBrPks131vPLFAeSQrACA750GWUXV+NfuQX3H9XtA2cMgip5
RGE0zH63B0wPq1++luh+bhowTQVRTeTlv/1QOerR2GJTq04TErvR/q2Uyi0Sf/zf7C8vkyZtRLdz
M45CSGjD+nNAf1fA5m6tnTGrsAGEZjTLitZ9irAv2/7DHGS1MY8UmwptoaRAkiu//GuOMKlpoYfl
9fAZKl9IB9XpIbWyjVo+TtnUH0CoMqznccWJzsavcP+fMbWIhCY1JBaBO5X88E3hUOv8ca59tN1z
X8HzhGYpb4G3hGzmAdit+oZZxTFvBOq3aTU8ieIkIlC+niIs3kBzh5RdGSAFtBII2eCK8Pdh9Vgu
4SlI10KE5SISq/YINni/r4KRtfH6NfFlGw8styYw4s4IMsVLSE2NZYTp2v4+R+2sGV/+H3nJlkZf
W1VNu3z8vEXK8GTnt35iTfIceqmx6xnVUBobkc6MYHnUPbe5GRT1Fa3Wis3Slxog4BmAyOyCAUrW
DX4bY0Njrd+c5qPKQKTZFiH9AzZpMaaBwSoAkfjXAkucCWgJ8Bs4dvSmAu6A+xA9Ho8iGRNaP5sd
1UkInhDSSXdjUJdKNFEd0n17JTBjZ4fsygPoUe4BZ/FVmeefon2y19GNQkhVoTRVhIY7qX3q9ClR
kwKH8hYCHFtcdhBgTKIZ9D4mZXqlI74xys+8WglajILFDDzdyw4Av7G5VtsR1v0AlMrrLDlKMMuG
h3q2QHd7MNEBaHQ1ZF28pJzcfKsmyJVSHmmFCtVvjDiOccPhOab0mvJvEzRJt/rynM27uKYdiqb5
CaDpFblULyWdRPZYT4daQzro/73Lx/xJt6tma8IdsaBXH/7h9JtjhwfGYXn+XmNRIAuB7V+u2lxf
mi7Wp7+S1BvR0/fTxO56jb7bHDmWQYHdfoZ7AZS3lDuwdW8P1/tqoFEEfUpnHWtnngUpCAMxEnKO
04FourZqxubFQ6TSjGq2INkT+t++21Byd/ttWSf5ayJxnMfVvV1lNYfpJSRpUmcXFDYpe0/cvTo+
Fzf1py0xj6b3LKF3lXG+pTOZ617+H1m1WX4jYHAx0Gj5eo69vLVvJo5F7tz2yfVAP6WTpnTgreVQ
cSj4+e3Ujo8qMxd2kVK8y+yDOVqzgtRvSDmir6VCJytqHf0AlCK0jUY+J0PFFnOMC0jxDyQvJ33f
kz4gNWWEfmFLKDGUAEV4OvTjJ+t/f93WjR4lU7Ul8jxISZAnblgIdkIIMJzaNC3LMu5px9PZK6YT
JJ9+yi+eRnAXDU/ZL2Yoe788/XzxPsmwWksKwOCwTHafUoOcTRKbJKCIO+PIKezU6kOQsqmATKsb
NV7j6GHf4RvW1CRs1BDghunesOqRP0pG3vzKdIxr+uTsr7xy30m3bgQdrbszjfvCW+J1PqhDDEjc
3gECTk19I7L9kvSqIsYkzYUFu0e9IMlKS/qMBmupC9EkWB1ocZAfvGpm16oXsomVGUy1E8VH3V1m
Ocf9pj3lH7CounMEuI4J1mycfmWMdqrFMOq01KY8LtVwPaLkIgTIbTtGXdcLpWkcVY4tMdZOVaJE
QDodG/J1efisXAX+Jle8RIpo+MeXQeIA11T+e5S2crkfCtHks+su8Ki1peRnqDOREWqY5SwFFzty
NZX9bvJxD5LzhXjzSASIIC2rdjv7zmZqYmeO5NUurx6aVkHAW8pEICBqp51YeuzDYjvuXz4tBJcQ
npzqzzXpXdYGr/bbaECnsLhU0OaiQ+1UPpscjXSIxzQK5gXNLTrLWMny6vUZxg5Bj3dbonSvDfOT
l25M4Y1pO6lvoGjw2ixzAnrOENph6EB6Lt4EjAJxIofyiluWXX8IS+N0s6gS9nCKjiDvwCLFPs3b
+4aS6BLxWlN6fSdXBPDML6hBq8BwmG7P+sMEF31SH2T4STqe1OA2LqzEdqOvV/AKT3r/uo2xHOgg
y23I5Guv5yPGXIz0+KbgF7TxaDa3zGsGtMEuwGptPIH1hRnLQ9EVl/ZT2UMtAcccjwHrTDRtWNbr
6wnJK3wMluHd4Optg3KGh6Oe6FQj4NKYnvHFF+Jpf9NLlabLWGDH/UaHqT5rqdZ385LM3BnJbUCZ
ZBTL6GplJsRGm3cE+H8vPxz/s6QfYWhoN+nCnPx2ZNvh2F8SkxXGaqdIFlj06c1IvZSVTet22Ua1
Poc3weoxUyWCT0tQ2R28JcRtw4lu7D+pLB589ghK39RRWON95ut+VcoYsdFhul/6et+Fv0Gp0SMQ
2wJ4YFmk7t1ciHRh8PwUK+GFX7FfN0J/O2ztJ8V83in1DKcR6QLHzpERhdJjptXipdQUZkS8c8xC
Ga5Dbzv0mGYNBQBKwkj4BsqpHtb/IeYNzDEvrdPTvqlw9+dcczRe2kBuuGOrPRrA33l18gR30mAH
ZMGsdspjYnxSTyq5TITHZBhWZhkzFqKT/fiiEZoDIa934sK9PjCQDRWIPBit5eUKQLy2fvTGcMvy
07IUS+XySh3oQVR0xXuAaptjcEzs3S7em461qb9LQxcRCcl3mpg1Oatf2NqsK6sJjAd4NFvgXQIj
r05+v8SXeidhpRSTQQFh/VBWxxy7q4kZlp1l8EiaaqjGEh1KGyTXLR6AuTN7YGTnE0uT8hPRuMAF
jd6I3b6pHArJpZSrv9BJVhIkjwUEe98O3bztE+f3E+Xicyq97F0daiaYwX4h+1hJ+EtZfebu9CFp
fu5Vhpxf05rr1ALc+CEenEeWjcXW5dzwVWLAFbAxx3AAyq0Gk5lK3k3lb3T9nmpBSzxVteOrSVfH
BaKSmOEMoHJ9FIuV5beXhJ4dg0zkJlvqsPo3B6yEXb48qDuihli0i92UacYCLZ3VvlvP+XF7TDK/
eFPFIvXPOT5y7VUy9SGeQYUKx77ihZtNE02nOoqHn9+Km07ZHJxX3DRaA8bDYNazIfqu0eMd7VAA
4kGDkCsl7EkGzRt+2Xx7cOZH3xwrN8ikLmgemyvGVHJP8mPoyEsyoLDcshRRElvy/y4RJl0Rhy3I
EsaLFQI24OVVp+5+AY6aSTqaed/++z5k+l2VO1YODyzygQ0Por5/rWoLT4qWhKMOF4INB9rgobtn
5VWQrPk4L7wIwhqC40FWcGcQuuViMkseJvaMV6emEpvFBokBgSgySF6GXBEWBdLO3Lb0C7S6DUdX
sloa+Idc+ALCKVgLbsDQeqr8vqMKlQ2WqoAtQIvehkrvxc+rXxYqdnK2GnyaQl0KcR9O6JVWVKbB
Qb2n3SsitVoEa+IG/Sw6/0JXEY+1kigXurjNTec5iyzoCLhbTBTpmXig2F1OgLN9qyz4yBwB3bQ2
zoiGav3XlmuBjsRPjRGsmdAuYoVdZag2KCbWnAydR0KbCHfw+/NmsPgv4Z5A+lPf+m8RoJopXqvR
VWcONzyiJR/E2Ru/YyLNJJJT3ntec0UJvJnd8QiaFuXZmYOBTMVdpn16o3fBfWuN16ybIjBdXD/v
ezQdeO+Bj7i9XTu6HW0D9FLXGU13pMlAJJnqLpDNRLr0cN5Z7pJtYhqDe5VT091HhjQE02PR43hR
gyYdeqVFeUzHD0WiuhP5OB4wcGJjfqchjsI8qEfKX82ekS/fhkucgKfUzCoxCtt+bYJmFaKUB1OG
Gs1kZrD+a44aYvQV3O9sTUzq/bLiovLih1ClUEfYKDkCB91uCpf2/rJQReKoY+yJ8g26ShZsSPge
a/fi3ngUKVDJkzCOGoGl5B1mnNMbBcg4vM0oV8It84HBk8OCl5k9rqJuFHZl9XtP+QNevlfZv5GT
do664T1AItjLZGrhQjFkR6HHGBfty7ARKSBFMePo4vDsjyvuswVXyLCQT3rx5Qk9SZOH0uDHx/eb
cIQAAQHlkMZ6EieVfqRcUkatRVQ6e3sji8QLFYJ/6UGIlzdNMvvMXs8ejHWsHyLjS0PcoSsPrz3B
UuuCqD2HyStTorO6teetZGURbJT7aTLTFDAI1IIcnDE+JrvKwcuWVwNpYLaSwe/WUvOX0jQtHGi7
oVGLhmu/l5li0puIGZNOXWBEgSb31MTTJfu/FT+NAKUx20u65Yl4nORkczItNGXARalYg4Y15mym
PhoIW/5dFU/uHogQ8VIgjjBvp5avZcH2GCuahV6vL16lur6OLzFG1fB4VPaENLExhwgWUAqyPhLb
i0gXAs45yLrIKhiTpb11zbvW98uQZSLXM/bSYjdnCyilM6Ny9BB6oaC10AkGD3FpKE2bCOzQxZUx
9PJhuUslnfadLLhNFezABhOcGYXKWZtSHrDeqq2hhzRbvI61op6LaAaVSRTpEBjZ3upi5WFKdTgh
05Wyu+wgXHWG8l238wy+hq1ilDZcgHpcmpWRz+2uC+3F77V71OSKrkBMkHBE2tt/z+B9gFTEP2A7
A01BjaIf6G5k903wdlGBLK4LpWxVoUeJGk3bVQiAZdg5XBgoQ87oDHEG1k7dmv1S2LlKsI8PpXbN
APbOC0BojNswiWyV5zzzrLyjLJppJO7K+Yziq8+Txyz2xh18wvkao+WvjyYLxyohy+bKqSKCX1Lk
USelccqWHnvO+ipRs5t4xBgnFc85059lI6TJIt2YmGJznoZinAZ7EKnVUNNgSOxZ4EiBaJD06PZp
Ee/57aq5LiKCK07PTw/yu1XadP4fFwpieW7Uhby37XQHW8w0SHbGefxcl/p2WvxbSkfcOEfCMyvH
GlSPpH6eTfTh1EvIYZsdROtZn2XyYwNwGfJZ/42+lw/yi85wVhgbJJL86TPIBNY/XSgdlcWrMX1N
NUx2i+uN18G9dZTw+sCz/17gg/9DnmEi6mXzkMfR2tg5D0IK2tkbaPADGezBeF0b+NkLW5T9lOLl
4uvU4A7tmezq1vKJTPJahkLZBKEf4LUNwZJYyFL3RIJNr0Sk3fgbi4iBOiL3v7icFUslTHvYod4X
ZH2fkJd3eRidJabCbo8oJbD5JAlgopPyC+ooHS7F03QqePbAzAhcYyAlifgYTCNaaoH8uVOL1yCM
Se3aqcWxdnbCIsCTXL8r+Wcz/Pqq0JxYrEa83M7QqoR53BtOjbQveFEBB9pvXwStBhpWPyJLjnl5
D2ciO7+CY4Erb6VPCBDJ0c7oQ5EcWV0jP5GFDgOA4ynDPTbT4CYC8flsU0uv+QRkHksCLQrO/8Xf
2v03vkRA6YOQR6JvbGkkqkSJF9RXM7vXh7qYrbIrRwaA8+q7gy1pzDOBM3jJ7z1xSlHAOnzAbOlN
etYal7VPQ5nCx8r2N9kRh08Hv+YpQiiq2G8yjq5ckbyNonA59F0rw6aIFaU0HRbgrrP5Oj4kFd2i
DC7LAZHmx1/CRicP5dgGbAEEAHFlxm/LI/PiczC3hdG+95WsI41KJuXrRtd4VYLt0P1RxBDiDegZ
ZV5pH/5blhXTZVAAjyv1Gg8e/F4VAs6Ahrniuhce04UtSgffnTrPzLuKg0V6+nWETYbCwTPA8HZ7
C04Af1jZGLTT4OhjFcGu2BMThl4zbEMqaKokcqy8cAMj6rBHoCCYG35BfFSwsXIFDOZJf/g+6YjT
RgdQVnnTlnWXiTAK4TxJaOuA5J5M3B8sAPyqTtUDxhDp4vyWqEMpLQE09QEkKM/fvJQE8xZCOC+T
MCw4omRfulFuR1I150Q10SBRjJhvCkhhmvFthRc4Gz7t/h3p5uXxbio2SdpNXyaQdb2UkKvvPj5T
U2arcGy8QD7OiyLIXxE8sq+jTQs4qNiOP2B+rj7d2s4hkdwo9PHFvvkH8FdzF1mmNFgKTfLGrPPa
tAmy8PWbVVDfNzKI658wmovABHo8F5OX2pRZHRLWO1x50G37SUF2jvpXAW9e1SmokBxcTcSJ/SFx
T7h50IshmNYTqeAeeFVlufCrNoHP2zDJ5XSmF5VYmQVt1F/cLlDMuimrB0MLEDxupSuXyTRAXEov
huSXP0f0SO3F7yd9YCOb+nGRbfJvi8KIjlFc3KAt43vrz1xkQItvU27o0KirT4J/sb5RsRa6xRTa
fVO/9prwwxJreRCp7HazapCyZN/nZ2ZaCcyZsnX71bWl/LjWEqOSYp9ZVQAMAoFeXDSt7ujsERWv
+XLjIdTZpbQBvzVSa0nv5QFVQRspygmg5BuUwQkrIt2hS/zQQuGt88dwzgdoAPEjeFwDxmus1+lh
1c5Dqx4OLuvJhjRm3hqAbUo+2N7q+Zls7LgWO8tSowrCtIOqYOaJWvaU/ijxHsOPLiVeTeV4Nh+J
I24oIqDdqwBEOl11FmHdasPEmk04fQ2DRQd5cnsdzcBB/YEFHChyotrFP6iecFWPqm8ddVdoEmop
wg+pCaZUYIDQ4C+gRMK9OKAZFyhazDx+HHl9ackqs6Vv1OBuJYecJL/WcBYaklF8UTghzUAnshB1
RC+PS8fzYRF3yUAbr6R9ShclYGa4W07kxXE3TTZAofxf6lp4OmfzntDwTUU5dhDfoLwHjYHoWiqM
rpBzQsSFNH3065B4KX20pcrjuR75CNCjS8ZPOOf1F6RR8NpAdKTGth9dUZ/GKPbKvPT1pRA2n0It
G93/R8PmMdNucMmYqFBA8L6nfEjPpXHzoa1OHsJc+8ZZPfaoFp7SuDcM6fESgh06AcicOA92M3M8
R8kJ9yLEwdm4+eLE+nEIXmZaFmTNWA6VaJzbi2maZlLnO55+QY28jdxTuNpzO9rkS5ncayAi8Mc6
7XQH+obI6cAGlpPp9TahzwNxG603tBwjrrofzs0228OULF9vsQSW3hp2LtY+UTmtdLHUlZef0Uor
7W/UsMEcGwr/Gq9L3GJoKBUGYRpLVk9bA3r9T6vYsv94sURZcFJ79CzgME2inJ2v/iplzF0+iwP+
WIdS7vlN6IVIDCm3N7XpfYY/nYOP3Bl3CbrMEfUZVhxqlW49dPLsAak7/auDEEWRWFQyjw7OH1gW
6vNxCMcYeNqJIQZhgHWqrplaj/5I16OhZ+DaesmyZ5DlIzeub0bl6SYLyCWH14UjDWG7NUCiU4x3
aG3+E74aYQn8YAxwdgtV4sYv49nuqjL/2DvdP0bFf6EBfiKqwx8jwmAXbtPF0ioblQwfu7QpFusC
5GMFsQRvDgFdicvDurDx6wn/DcuAUxf9XfXdEX/qoPblNdFvAheiGqsIPoO9TsNYwbn50YiTmv/0
kCPbBVtm9Y4UxqtrhFLpXMCwTOBbrl3E76SBdY/O3SAffupRpDUl45LUMfylDodutS4dPoZaO/zq
LMaqBJZYvQKQo6xzxZah8/brBDCH0GV/u1D6Fl/AW/KSYch4osGLG80hP6XbTenq3fQ5Mjs3v42d
84RRQC6IolxEgvztp79qF+HIcR+P3qPClverzQSdQZPjNt99Pj6K4h8K27R39mgd+FhAzRY2VitS
mOEoxBPMMvXCzTpUTRqDDl2wOMV90tDt8fykXyzhqoz5s8tULiSA/RTND8TUElSuWDPsbdFYRz5p
q4g+r+JcNWrjJ+aeEv9atIowjXYso/4howtLJldTcjfDGsMea/uiIWawEIyg5Iyj0rmjVqsp23gK
WTtjJE6l7DYcMzlSA62kUQa+ahcviceSWNtP+9SRBCSS6Se1IumbFga2WST8MWtQfQyNpPbjlR/E
ys/FoAVr7iShyqGXHtWKtw40y7V0ry5VxthalmD8/HQYOYgYJAD8PsJ0vwT1vsP4mnJsiDYxvHaY
x+LQsJBfoytrncXv19QYdGZMnHOv3GIbLZKo8fCUHxK4YrZRcfg2J92cRQH3SivtdvB7MDstQRN1
hxnJLD47LiynxDoq21sc4qswp+7P5wdVo47Hlv5W7PAPE2WHg7V99pVpjXQt6/HYYWCbIx6D2OkS
ombr5P52adVgp7pNBc28EIuc9P74wlPS+wCHAu/4Ny2D0JTMhzq+EJ3LLBvbLP4vaVpGLbQYK7uk
3Bj6yn3yMMufv10HhXIEaaMsVwCMf3BvrudUhNQckB+FjD1OGkQXkB7zJccPthh0h+08C83+RWN9
izHq8kDVaLSpUjnxBllYyxRpmn0ugkXzMpkydQPFqqlhSr8lpyGSpKnsK0LE2O1FnbpYw9dVafJj
N5IFX2k9eY54u+u/grDBVAwY50ivYt7/j21RwVIjkq/UPvY31vutLP3aDjrZ4tHGavM6aR4Br5t2
9YgSZAq8CdwIuPA/bKBe9k7rg4FByVEDzuW3c+lUT9v//BcNhNcLIFuxcDf7PUMq9UMxm+IxmDqS
MbvFS4nPBMCiE77/Ps2hUEUFiB5VLIIQrcuCSYMIZu89BAh5sixnZjRGd3riAj5+DUp46ESnAm2s
NasNSUUCWLq5zd/PJQuroBOM9HDnRid6KrqsrItz27RW9+tBVG6nkCe3O812iqlawB3jtIttTmdM
bkAbJnggQdQqdGGFIhfSw8qjhRC+qI8Agc0Ldl4Ucr8AsHQfa+T1fZ4MDLkUPtxmD/bFTO5/TO1r
U+W4fzqlc9rV5l62YudBbaea2O1wlIbD308iYgnPDc0/s6jXeSPGt04NGlEiHQNfT5Lm6ZDyayBn
eHZ1tfWDhAIm48g4BJu4VuO8+SREGNlTF7KdF95GisX4NWAxxNfjIFhvicGostvbZJrE9kpZ1y/m
YcYczyK4J//lC12JoHRXKDG+4cq8Wz44WBWL9n5e2bzfy4f/XtRUXdDX/nkax4d/AFeOH0tVByL5
ztgQettC1tUJLSWi7Zn/1bi5BPq7i70lIWh04AjpmFkrvuza3u+tcleKb31ELbwCYnF4aQcWdWX/
fw0DtQjZEG1rSMYPHi3yltDw7zikZj70AigrAT3nGesKWg7rvbJ7rbVicehis9YmkT7qBbj6wcip
8872UCjY0OAn800BJHoGZxDdZrP8GJ+WxRsHo/0kGjbbShqeG1fYONYamdAb+VcWHhfMe8v8dbJp
4F5quFBxd0C2MiTsyY5he8GF7qY+XaEy1vcKNeHg4R27wI4vQKC411uaj9fNo54ZZg+2ITS4DCyB
VjR8W/hhdnT5cfcDHVxkfkpxdOY+0tPVDcUAz7DDM6MF9CFRWi7lrvu9YA3PU9GuwBUTAb9/OEXd
3f4vwrf+AjDan22Zcud3EiSY3L1+hZbBL23FnkD4KzVU1kYYN3oqcx58HgY9n7d2A81VdRuy5HG7
k/YWmEzUP3c1SSMh4qYNirjQh4zufpKTc7yEj6XkP5WwcZcomnuaF582jKsfxULcV2LoUgl3ODMu
I/qTCzqBKL1hvepVsFByKyxrTMNxvFki8W0NUEVB/zuF/MQ16vVn73QXyMK0+d1y4tam72iNpNfX
OPCRLtDeMHWXLVPZi+qm7jsjY8MNVNBug+HcFvlzCuUXhBiC8zQbd7pC3eBQfii88r9b4+1VUilC
yKqEPqLQrD0vZBXQmENbFVa5n8p1deJ7Qzj8CYJXYNsE2NDKn9JbUN/BkQjJqWg2iZPTaUM8ssmY
MaLpsY4/tNq+vczEj8WOK/EDnXC2vk1e/oc/LFHXbRszRITaAkMbMphCwLbdntX8wafbkynG5/dW
Wn/tAMgc/wlUbfICwje71H7ESqBGOTNRQQHALg39eGshs9Ly6hPRT7ejy5RZ6esiM3HA0ekxdVAa
8oJS6JF8xWPJBQmC8r7nac5NdoYxOgN46SbCPc29CuDj65fxlrC8rRmpqpg2+yZnxaLwAKseTEw7
MP0oudJhkxZwfaXXDC7ieUyxkTh9yovWO8Q9t6a9ADPik4aD+MtQFIQAWB6OlYJrr0+VVW1n7DjJ
j1ltbHzIUnD/C2MqG7sJk91kDcUkNSgw41bHqN3TDmImxPOF12dASUanvb19lDPx9HDk+B0BY+0O
Z/UF/Ug8N1wiG2Lo2BzoEXBEYHCVQkaS+o23bjYQUnlBTeAGvZhoAk5GmmZz6JMHwgU0JN1beRXg
kZq7y5ZbwhdXGQEbydj4tLTStdSIB3pyzsanIkwC0xElhDQyWfK2DUNkOA9LFnzsLZBuhh75cXwM
SNGf3zI4/mzd/OB5UbsqEP95ytDve01ffRKoGTCylGL118SsTS2slSJ6O3qqXK8fkqy39IUYfkS3
+oIdM6NUFZtk2J1+eGk1b6KoJJBS9LhrVEIUfV8LiYq7BSq3H0Fu4ePtINme9As68us6XManhBO4
nHg72u3ZbGGmEgmeo8HcnG1hRsL6iDX2IMoCKkn51NNJtQe6s5wx+sHV2QyfYZbKm62c0Xpmop/U
sJoOjaJekfaAS0y78CFxQuB9TVEqe9JaAErft6RZ1mQCdyv9Z/w9UeUVru5VGPpQNZc6Gkn+wMfG
jXLzs3h0zfnEj0TD5ms1SCvJRB713fEUOdYpkyJYcIzf71JJEkelr6i+Zi/Pk+QJRWPegPDRbjxf
VQ2mjXP5naWNW/1dfJoWbjeU1HuD4XSNd15QUSZHQKP8PzQaUbO6voNV9eiXqP4KKEIw7DGm1MNm
h+yDKwPG6PVPpKQ6+FRTd/QAvc2wA87RTOMRLDSuTjuqVe3lpYyDNT6G5IcrPdjrIiVY8890XGLg
YYorzm/HdxugrDNwjS28L5PYtgsK2xdxOXnrEdg5jdFSTc4G3wpH1no2Y/VFo6aaPDSgH0H29uLG
FrseY2n1IL8LVTW0CXjGS0qIYSTMRs9PWcwZNYPOxFIWPuwloUx3FRCaLP8RlIvpquL+L/NOABLE
TbR4U05JTKVuGJotMQejkU8CPadwd9zU4pNFZIhqT9x3NLKkntIYLFZiv2Eg1H7CmY43nh+ReSsi
sGJQOPUToFUJLX+klxZnL+nUO7mvAaFXvqPuoK2WmmpuGw7P9MAXe4l6Ofju8D4elU21hijIcnSu
cyLwmR38plpH1aVjH2rogQj7lHyjxkmByrOh4XVaRg77FyfQGPtkcaEx07YKrCA3WA3QN0tnhBiW
CBhEyL7Db+CjwTLS4F8ZGf6UeX25oRDW905D9vek9q5mUtyBiw45jLZ0kTOk7LAMI6tZfG8+tBCN
WJxE0DHDOjMa75c/i8m7vvvDHhzCH56SymzBTZzWnyhAPH/V8oYhyl8hQgWxFzV/F56kS9/j0U0f
FxfaI6n81h6MpVX1ELoBJWcBoYAzTXrceHmtOq58b+Hh+nsPoCQow3/yA0xrjJF5aitaOoqa2Teo
EWSO1xxIJfkoIwlJr/LFDV3eaNVO5yXvPQhiY55GEfLAbdnSmTt75vLlv6zCmTFZxyto6WFr1V9o
pTi8hMXX/ZdX5yFf3mVMoLbVNQajbhqPzAGesIovVy/mCqP554PdqEggM/7QwA0Wc+pPSw0JPi9C
A0WPT/TkORLsu4sC6Ge7F+at/cB3VLB+YYQVyZmms6sdeeVrtLLxOMVsbXmeWYiLe5WjEbv668IS
eTz8yhdO0q03If1zkMkPA9sk3mLIEs0EVGd2rEUnQ8h9JjV6azijkC88MZ1QMOM3YAlZIGwLo6Mf
PB7OMbnWpT9Cvl7YpPVHB8V1ieZ8qWJ5TUSV4z4ifhe+KbNPV8Ix07bjgK/rJT7o79LBBBvjrT8V
m0uVqLf7wUoetLE1EFtk6s+2uEmr3aqiolBP1aM4cDIL1RsTQ3XSOH/kZoxktbMiTC5g7FLbNhDB
cM4BwEYEB4nXtmwlyV6d6cyPsCdjXzP9QsMLQqC29KYL9yG5EkYnnjSluSDwDG2c3ySY73bdRcGO
nvTl24f2S0kCQwVFIXWMnQjZVS6W15IQxcH3MGs26EieIkHnTD0TpoicdIzFkg5ow91kRBG+28vG
LkAtZnu01Gbw7Il2BczspI2CrrBsuHrbEQ0toCYOb0L5MAzkO84FDowQaLjD5pcqeGCDMIbTExkd
XdLfqDQw8rIqfbzHfioMX1vvZJwOGgMxBD9GOhuYOj2IVJuzMOOvJf+43vb6ifujxJoqpfu7DC0n
2yDDd299D4EMdVnxNHPB9vpZWNkoNmo85q1JGl1FSbvUdSZDm97i8uIgb+XvtqCC9LsBl6e+Gw8U
d6uvvmLIo2lb4qIXQMpQac42HBnUSLayP1z5oIBwBryaWhLhnWJXgwzBRqslso/OeCK00GORsQ7x
/c0jDsVtSc0TBSx7R7UAL/zNcJDwVGLbOamljv4xlIcUOTWzdcTm+vfUprKoFZzUpFF7320SmVLY
tpecK54UciCFwm7fBW0wJuUTxVU0A6MEb4fo4HTJxE2k5cLNlXF7HWmgiXExMt9DEnLqhL4foqSn
RSA35Z4dT9AOrbeEpgIRTaGCZWKdmKPsVLIL/U1qPgxSAdH0lmK3VjlYASfonIi5/8MJX8FfNwxl
VkH5QWbUxvIigOlMYOAw2G0mkcOcMnmPGkk9Ze+UX8chREYjaXTONAT6oGGZO4RqJsvVEjAscsN0
hHdNV5bSKatQeVuzA8VaOB3lISawbMZ6du3lou9kQoEYCerM3Ra5ArVc3uOggAJeWn5bvErtTjPe
4vGV0b9N/NzzBP5ERi2P+wZpRMaOafrWTR1W6QcpWiu8dzA/QGkWsjBb6fm38vSxx7ZQtIbCR93E
o4DYmsDjIGToMMUyWDCk0/VwYCZx9mNrAyDAJnZwZfSRET4pDw6YNtQF5ziKiORhGD6kRbcsPGf5
CRfRGrnWJB7aUjJpXuKIEfgnuX8Da2zGpUwniw1N3LX7Fa8HVgGSary7OuE8/5YToCcBJBxuLsCW
thI/Nwg+4UTuSq1UsMicY3Tc9HKuON8fMBlUXMlCdP8XIAoTX89Q1ir22lCwucAAetpmroXSUBud
rb7NnLPcm9WP8drX64bKf8C4KFBHz/aR8RHOdggvbv9GlN5g6KY7KQgiqbiaCj8XYP5laI1Qk6ig
7OAiS/+mRQ2Z6+YKPhS7FeHFzWDB6IvR59A2fKbZvJPgwzbEj9Ofq2kW9AevXoHgkpU0NB/dVS1+
29dB1RHTxqDsOf+e2pmHteHP+hVr8NDE4LfcEVgTGxHs8tWUaNBOhasCbXDnmq7KWjDsrQnY6+et
cxchr6W/uj5e4sNKDd738hqYFCqWNf3IWoGac+fbDCBnO4N4YYZ5P5gFu7HpelljygjL+kiJLkER
W+N7UFi8917RrZZXxlAijEfy6AXUpwOe8ocbkMtzLLoYTIrbAZB5xaizNK9S4hn9p4I5y3MvciOL
3WnBQKXgHafARMbN2D8j5X+DpmLaWJjwybLX8cvWKqwtcVW19fm7o6N9G2rw+irbm3Ar8MM884Pp
akF+MEKrzJaKT8OodnPaddgh7DjmRskXghkDHvUY7ZgYnxkZTxQSUjfkqZb079Y6P61gj2x98+bO
LHO/IECUMzcHVUblu5muB7FPE8av6muYysui4jVVQ3AqrDZP40FtjQ1syJFqkmF1TPk7SspNyH2Q
0awUcUX+/ta0sJIfL/XIhKru3WG1flqzRXwKQvGXOKI4D1borEkqjw6LoV+Ct2PmAuFZbcOtbQl3
sMIpnqO6NpoA4M0Yv3sciKsuixZ+YJdsOtIyzYcUCZCvj3U0dq06z4VAs3PY9/2agLU0aDmxn0oL
532AjkKeoj6dp0PknuEZYewj9sf1ZbIzR/6B+k/y+bR2iZzXFb5qhspvoGg4uBfe2BFMDQ21mBqL
MAszjbOeVd/zjRblcBiFr3SGM44pFEwClMv2V2+dA3Khz41Dz58KUJ7QIAzgcYI8IlLBGlCbmhnu
FxmqZUni7HhuqGbJuOJfDJibhbqudhDaMyXG9dv/555FKe+EuWm1xeqY1ar2jNrdkop3F3Mo1i0p
0CgEgSKQMv0U0U2fnMo/jy7E5f7D8w4tt9CeXjOMp5wD7a+QYjyrEVskk8h8CkA+9nXy8bi+bRoJ
7XON5JDH4COJtf2Y3dFdNHLoz/w3vAWeuq1wYM/IZ3srGX6Gtj5AzkHpSRFnkxoaX0klmR2wKIof
qxSPRLeddTeMeet4SLoMChVFuV+IaO64ptMwTJ7ubuxJgQDw+W+rKzt5eQUr14tLsOuQ3KSTonFS
EX2HShTpXVjioV3alEpLiyj3fp8R3AOZ3sXEPbzan0uUmuJi8ObTLq4s6IHjk/q2JkMUFupdPcv5
hp4uEvbEz9YTona8lQ9ZwPKcn+PN7eUZwklg7Ul5lB4R/1Oz2AAoqKPFMFCwJH2JynTisFv/RQi2
QiQUCLi7iIIscR32vrTqPZBqHX3BrjSvoqBLcrsmHAjV1IyiCXMFiPxKyXRIqgR9YaguJjWreQmS
UAcCGCA/YrUcwTs0snyEq82Box/rQgp3u1rmrbZIihra5RFAzwskpUX1FB399v64ibNmTfl6MNfx
a2TAN2/Atrn0efIfvF0iMiWfJ58RDvTZslQ2dZf3atgw/AOPJMuAPFiL+bC3c7GtzTBtuODCIfCi
f5ya4PqbOyIiXX95AeQ8SMVWl6qKRbKbCG35ES4F4Nj2EMDWOBSgS7C3hPPKPm5YTV5flWR+5jPx
qTdHgSX2ez/NwN4JYtzAhtafiPVXcTknFU8x65dRA4C8wP2jsFkoEWR46k2EC10bX6VV5fG0BGOG
r/I+bFil8/YIUOTEJqVevA0GGTre7uVy1iqL1PZPqQZOIAT36pucfEbEpzA6PL/w3uyNc8RJHQ8H
Gy9CoHk3eWKsVpgnuBt/Nd2okvJxF05iy3agj3mEW3YPzTlzC56vc/mi0jLdW2T5x+NulrkY4me2
bWXfYYEqZUL3i8jvsBsnR+vSlb396sFdoFO2fRDTVM9LfW02nZOg1IhO/aJWjBQNESC791+Mv28v
cc1M9QC4zHUsCBZSQKyZqQTZDjhiA6GHlm3ydzGwpgc0ee564Y3vl9X4rfhbmvB1nbFScJ/6k05G
Ewo3dn0aeR7qKxVfqw2Ioee5Lhye7NWHFm/f+N5skBlC3kiI2mN1bIKcLkdy1EZqAfOV4GzlZ7l8
pBqqeDcTd9tAQyb0XAWIkH2wP2PCQ9k4mQtUDqTsK1SD5UeZznW9vAx41ICclKBIlv/Th6JVyxp1
h52GPCCvMwh16IEE6yK7OukQPThZWyS5X98ZKe8qicO/nat57ecK340rC0VqtFFgwX7AEnVsi4Rz
F3hQ3WjEWnA7mVskss/ixaJEDgTRIx3PL/SjcdQoo6k2VMEWA/w+aVemMceYU4qNs0LPz9CXOSVM
ID+adXjIEm1bE6Mbz2XoE+oO2LdmxS1qDDZyvS28WYyKTGVgFhWGhv3GoZUUMEDPi3DBEsP79i5x
47KKnBs0HIrk5mC1mW8ZUn5nMj4eCfJ6QQKD5e/j5vN8hobPvVrqq0KJgQ1G1h+EG0ReTWVSFCWy
JfY8HGN7t4fQwCK8ADORAvSPpoWTlO7yigTCuPytbgwcFJZ14he49bQgnKaLqroY1i8Z+eZIZBKd
QRed1dQ/KOriz3QAQT5nKofShXw9l2bG8VtC9ITx7uqjXwSbFJvQAZpVv3oiFybzSY8e1aOVbewA
zfY5Q2WIYfhxvj0XA7bln4XdN8bZ9OksjdWa1JmLjqJ2boS2+c5CPWpzuH61AErtCJ4DTPj4Qn4k
GCXMCyVK58I1zn843luovyWcGCgzCGCwx8iwjksQ+5ADNCIoCIUazop7EOSVsP0benSwn/U7V9Ad
b/FvsXG77+nceJd4RwOH1UJQ+Q5zQDAkp1qf1oi23mGNnT1OE5MrKRXdQsAkavY+28rMqrT6b1Ov
/BV4/PYGBuhMr5wj4+2nwSZPqo9TlB4oNxShes6DKZ1qCL77gGT0rypSV5sstXk56g8HNxFaM5up
GciaXDoCEuBGWagrDJQvz2C3ZvCZq5iSO/scr6kiUNlMrAXkEAQ5UfUOVsNYVfiK7tO7lDQA/tcL
npJu7sOUI+qZDSyy5aIJ8aYvu+U/7+6JeDaiYU+VJPKioJdFU2WOt4uvOij1+RmOKnh4EXjKcW6P
fUH5EHH6b5m+RsdSKXJB6erHLLyxhrk75E1OO+EF1sAyQ7/OgZQxcd4ZOnMtgRErgthToDCuXMsI
sJZ866lWvuGfEp/vS/0w3lMiHGBgZezpQon+3wW1cKzg1cAwC0gZhddnm5TUGExSidCRv2XdA1Tx
FZLpWM4BEh9OMFfX2UU+ahwHoGl5z9sYUZNpEl8aVnXI+hGAnmQT/nPSj1CUWh504Bx00wXKNxQj
zUaNK4te++gNj1qtzA/rCVH6F7EmjGmdscaxN5Jy8BOKyOy3WwgJ71zzwz0wI6yks9vpe/O9m+1w
xmm4KakwzfaqVlcD/vrUokri+n6RUqBRNTjc2HPTd4vgJaKV2ow4xs/1Fr0oatziKCmPKMGu4SKO
Lskxp+/lzHTam+EBKPLfQfdSwurIV7X2fi2VWuIBZ7iZD1Z0xk91HAeplwQErVPx4QIfuf0WQvjR
uinXQn1a94zg3QMIK/97XjDoLLTa2cw5aD/1mnsPyJD9HBoov9wTXDMK9/wrVcArCvKEPrw6IRZh
d/NFKc1BxU7UeFZlkRSmXLodLVqIagQLpsEg7hcc5aqKImzPxmVUul/INk9h9LoC+UY8sWpzphvx
+AfWWnF1rDcswDRpC1t/lYXyQUa+RVw2SfaXKwGSumhBqZRnRV7AEQRbHNUuY0R3iz3ssMOeh9PR
8GNybutUCsiihhLtQhHBEKfvShDMQVhwxI9tqu+e1dkF+GYmp+sor4plGvbK2qNABRACjMt9fcqV
SuGtmP0zQeiOWILo9/y+DEITKSJGNirVI2KtfOStarW0fkqo0uLUq61erxRJtDNww+39N1uh9g2Q
EK9QVa8SG2hI6kL69GYNAFn8iGTDRl6ym5LXsOZHeglsHm7ws+GuxnCUP0w2JQ5caj1DK3ovxXWW
HvQ+LFUW1/wmPf5AXpzCjaqIhisPq/kpf/N4iDDMSSKLTZYnYkNITObkBXuEX6UyXTA4INyL8Ryb
WnHXWbbJfu/a030gsFWnGtn9s8HdDz4e/0fjDL8QX8KKRmiCuf1LY2ISh+83e8j6aYZ7AV8im0Qy
XNx7PkNgMsf7sqes6KosLDHV7a5/cme2XJmB2S6FOtVGJuWBrHy+9TBS+yZ5YbqChwZFKuGGgBiN
M8qaVKsNTRXY6xXU8IjxUuXQcF0GCY8TF9ui41FomlKop9vZZlneXmN8e9e8nIAqHIHVmCmgqlHf
DlfF74jRrEO9FhprYnsZEwCqpnXSv/huyH94L37j3sHFpOSxgcAyHKb5FE7Ss5UfLWQD0PxnP0ji
/+Vxuy4IvVAu8C8O73PTeZtbWqMGDN3wxiIoooCh31/gNbTgCxT2xJ+Pjh94MaBhHpt+dxxwDrOH
elfcLVeP7trWQO4D6JLcq8XwyI+ryH/91Xaw/hFy3vMymlyOcYMCEdtj2oSaXXHjUlLaR0/Etl/J
NEYu5mZXLtITHNdutjcquBUu0oxnHEDEXJyaJu6QfaVNM1Qn209PsrMSzN4OG5XLq6QRAIYSmpXS
H6ZiO/8SDe9QOqgZeRyIibYgL4OOakRiQYakFyS28a5R5i/teRXKE6L/uiBjWSlCM3BHGqaEYJ9R
R6gns42eoWpJyk2/KF76MeEBtuxPwoAhB3YMZAgXPlrNa63K0q/ZzweUd+7YB8bGcz4W29ekRCYd
l9Kgi7sKRJ0U7ZGtir/gM82WNoBq8OVUeZDU3QqPW55UCLhYqsBhirlFAmG1+XapGTmHdn7A+J5c
bzqdtFTQunswvNiKiOpf+bl2FTEl5lo3SsEkG99ZKEZpwRmgdOom4CXqBBV/smTcNiN8cB1Ca8hB
bTSM2m/uSTbNkmHxs5kePEYr/nlEqvk87DzTxfUacj1by+e/xYPECjBVjcqo9zf3IvnT59f5sFu9
el30OrJbNx5CU52L+Vw82MZEdizUSXNxs9DkKBEXQDNqrqC7uApWMFk8XeX6LayprivJQog3y22m
eTCWJV/yotx/bZtJJzsTjh/dL/S/tjoNz8a1OGqhwCeHvX0FveqXQrNV3zJ1v+rtWw0lvbnH2mdn
Rl9s2ofepoKG12EuT05q7Hx0cs/RWH8430NtA5k3mLxf3EqZo4t0Qw+CAgxKjCEjZ2BziRkbdHkS
DrP2AXy3VRnaycfP825r9w8d2T1B+rPgGMfA927U2NRdJaROEXAU+wUFK4otu/amLPRmZ3T9cGUF
fIagwRyAftYJGLh6gaXXseZSWRwePwHJl2637LR4BUiHz6zywgo2U3MH3+zG0tY1aflmw8337dvW
ES8lgDlUgN6Abp4OQBU5J8FoPF8wl4sfK7JQyzW4r3nOeM+3soop3OQvu24FK2lBSx+dOK7YH4kk
ymdCs7Unjx2Tqa/1PtsvbOCKuhnqDteLjkFhq2/CWcdS/ed7kv7LJIvazbD3oRee1WJkrQFNRGnl
oui8rOGHHPEov/9zKA1A0/xnO+2B0GpK8ZfSMWrKT58V1Bbg1uQXwp7BFjAppYjXmlKHoehsrk7j
ZIfgnmMslTQEu45Vko8w6OBf8amxUWursk10BcrXhnMs5Jq9Wo/vMXSeSjlnm9RhKiLl7ttoqNDM
kdc+Qw2r174BDFKA3bTL8FCZPzmuDzeYxY1V3rbwmZBjsONrxjk1N4eOf1sVlRmeXMXppJel/tf8
1GNT2RxG584jFvV8NHWR5JREG5V7yZCU5z4gABSxEjgRvhK8ofOAjJOFbgGeIQEOuvuRcX7alWG7
jVEfswvwsO2yKe8tOZsqdNUerDIxsfeZBTyRiRklJ/0adty1Hfv4jWio0Z0YAN+KS3/0obW9DGGR
vAvGxxNo1llMT9TDjf5xyvC6fS1QxGUDKArdP0AtfenereLsT2kARoZ9DsEzibmFb+zt7Ir3ywsu
BhC0c4zca1VKZiDXSTukRd6itBVLAEk/En9/3VcYZbssYE7WVkF6o6qYrrA//ysOng8mdl2DnI3M
2S3guOjmbCiW/39hDyjknUOPcOeGb+IdxxJzsit3qg3ifoI+8B4BXwq9K4whQclfqDqrJCDix0Lo
Y8/rtmBykmHGGr1jGs7bf+FtfW7t8EhnHc1kMjh/HkP/JROPJzzx3M2EsEwURUMzfAGYhedHk92C
83AFo4D1DjxbJSaN7E5lAaH5Y90QHp5buiZkaHjKh9aJ5jFVi1lnJJEXxVsuZrHAjLRALgGrCfYD
LFAux0DLJ5+Uaja+TZd0XT9evvPYpfNMSYxHUdo4VI7vim1wTAY4xhpL4f86fS5QqWtMnb6Ay6kN
4Q8NFS5Ewxi4lHU9RIpyqolqwMOWtg0tToU467/baxLxNPpSeAhRwLEdLEqZcHCbqn/AAbYxoMkD
YlmfFMbxBWEGt4t0a+YXQdL/lv7br9uq9M9spz9lWVvGxn/UkqA3lqhT/U6mOsJdyTTlQ0kg1KUk
ZhhRv/EB7T4oNWiGp6b3tSzCG3dkHBGlSS3mE8Moid7DhL85Nc+P2hHl1qCYhyvEIa492RcrGBp9
W9CR4tmrYfi9Zuj2E0oZ4me+rTdU1kGy6vjPET1SdW9JlrklB13qvjEAcRasxmIHfGiaZC9KM7T6
jghNn5iNQ5a5swuV+wxLnmIKaEU+vhj/0dvFQHNK7j81WyBYXq9Oc+GU1gZFlNEY2XAmS0BHwAQG
tKW4rhQCuzStKxPBLOARPwqg+JvFpWaMp6tX/rBnl1iSXkasL95RYYuS41n7ZeikBDJP/qG8V6r3
LhrpAmRhNHpTHC+054f9GbQhs8tJdw1sQRfG8dO6DDYQ/KYxTCD9SL2li/o1ZI6/8aVBI3kpYCJV
3xa1gp2/8eOAnRVIwCnYFWmkeIWgEFH/y2p4l6VnHUEHOzHuyqFsPW5JIuHnHxrMM2MOdrRZcTXy
Zw+340W2WE4LdeIg0mrRZ+wE7uWdTTE/bXUnipIQkjGw+2UA+8Tigh0ykTGe4/+LBNIsipyeNi2A
IkEnVxE6L+l4qxdxW3QJJ8D3rRPF6QRAEJazx50D57Ej1yBBAlSvPhuavYQWTKV2CfloP9txoacm
6li/guQJUPXWVtfU/jWThI8cg/ToC+HUMves5F/4patLEc6qheqhvmpbvTU8TZTJ/pDJnr9May1E
ZYLFIipbr5wNjsrOR0jlZNinPhPqRPy2t0aw0NzcVGTC0/13wMqW7T6iLwP6QA1SYvSS3DzHso93
Gy5l4twTs8a+kPoEEjz/Q4eTnikXEuaL29r5nP+fTmwm1LmCfMGagHzPuSqxjo/s9CkpzNGrfddq
aMWABFhOotQiymcfgfJhyJtc85Jg67yRtDmQ4Yz1Z28l9d/u4K8AXhmVoR8kI3CzlyMB1NumfrLY
psV3rwXvl7A9FMOnCkIBcwfWJQejyleeReMfAGrS9uqQgx5H/H0OjzDvJhe4dc9gCTTdbT2OO2Hy
1BLrjeTlOcdYuymO0JO16NffkAlOT/atG23FcUyvf/0LmGDMQhJhjEWREUhAhzCjMWOidi9hp26A
PDI/DYjRYj1dHLTxBfqUd4c2tTtMInez62qIc0Y47nrBRHWPRBVxe1y2IqB+1oKgKFpcpUD0TzX2
5/BIxX6VxMzyuevTu6kua+R1Nkm7GkD6J22DAGNRVOMQCUGnfZLUaFIvKP+yBCy7EqpaAka/eALk
KBxIGHfTLfAfIiQ9b8rgcLTqWECTxpRai/vdMhadPVRTIEYlxNX3tboAGSbbVa+RxWtvDKh9EWg2
+qL1OCRCJRzJ0qusoXLB2T5XorAYSSUWxOpsLQLC8obMr7QnO/R0x/1ndIt/4dG7ndszzwqMqoiN
aHhmMIzMnaXep2C74ohmL3g1naRtKGJDj0i+SsKwhcaz919Jpv8KSxQtLWdNXebqO7mn+6ombecA
OYTaI+G6j4bwZLyii2OqHjCSsa4yTMyuG+5ONHquWJHwJitengLDAyjdytynz71dNsrlQJSdM8hr
kRClw+uUM3s9s6UwM+mzXCW9PWvafY69gvU5S1uimqxnX88wbLMBaq2InUjlEDiXzCLedSFeC/gF
1Zl9jdlprQanr0LdRnLE/WBzCAwEMQDPb0qgKFxpUOPD9tJtjez/nQPJ4S0MknozMAwZBeuZ8T/x
F0YKophari2muaRhgqUA8Ih5UYj8qLUCqYuha+nzQw4gtVFslBctPe6GeD0gzzBBNCuCtCA/Ebyk
KvTW57tW4d77tixVXqSmysZ9MgCxLEuRed3aD2iexPQfdrj/VZtImPMFbCv7qTTohJujFyBkLBJh
lThqvfe0jF/csxiIjc2MlX5+gLxxqaiND0nKCSxMwye/9ek0V7awg8sow5hEgRuj6Q8ioH2vRgJe
yV9b3aaXUftxuUAbknuOaN8ugBurZzRuLfsx9oyKB1jea/tXWth7jk+13HYvw0nPrPT9rAWILR9u
WuKOUMHhG/RUgeboXgxLerqUYfXvswc689oZQLNGTQpUoNOh2dqPMRZNIjkV+ov8E428R+HKt1yB
pBApUZ4yNAUWyDdq7SMmmT2au86FDvrAWcUpOc/6W6ZuAJrB+gnplVnH6jSONLdD+s2zufmAxCVr
mW6C3FBGUCR97WXkGLVtxOXUKs20ToBSbV0cOX0rR5JzRxUaCF0lQv1LNog+eWuu/KpM3blg/eo5
ycHSYuTCghos32g3P0HGMyNWs0IX4WLnNX1Ok5/aApuUPWJzfRHOiUNRxiy+61ofTnNTKHtYd0uD
gylVr1h1xPy5GE+b5rzTUc5ZZGChgsryy2KBXjHgOuSBMRl6ul8HZFfGEDr0F5NfujcW5o9FzkOC
nxyzxpqA+/KDkTcr8mnDKSCk7rCPFjQ/rDFBjCO1zv9vMIHQdUtmzIjC1j0c02fnBYx/nIR9D0u+
e5/BrBGLxlPb5cPuOf2pfVBCdOID0UxBKhYYKO8UdZ5/6uj0J08PAEe088Wy1KYfQCZm1cb0Sv8o
ksTLtQdVqNtdCO5XW41MMo6BtJdWo3jevuGGcCpxoxfdyBQg/mv9Si+bss+oenywp3BmaqKi0Z4T
QgHErj7IU3MprbU5eG3q7t4T2YzKLv8WhwXePxgrLFhrlSzi3LMlkfOIcxwibRK8Cd9htvm/DV2f
mY54iflAl7s1+dx2JRTeHSegnHhPg4THqluTaKIRtEGG3964UP892I9J1iE729H7T7k/phiPi/VV
5UPyflZaZE9vmS8QRvrg/ce5TpdSoMYfp2YBrDFYlbwn+jXT4BMFYZdYCfrZijelvdE9o3/dJxPP
r6k1Y1r5xAVSTEFLxdYYOzYSKhGiU3c7agWzUDQ37qV3OGukDjSG/tgLBKooU3SOjsadEKWlQqPI
2rB2lDHqPxksktuNJhZEvllkDxbW6zQx1R3yPwSrvXiyTN9Qf8HCRHUcqusiXJl099bKF1l9h5Gk
sz7Gy+HOcpfHtbrtHsWGYuzMRk1WAaBcndPmP7hsNgJlvSMs5ls1crnQlpye4+aduiMWc677dooi
ccodRDGRrMITQ+bXdF2vJxtvvv9DHfjsIKYWze/saF6+faKb0v/APvYJNIR90AzRaXE+gC+eDmdh
cqYugLmj+3p6b7pJFKqkFcYtKEcNYWi7SggbMXq446QbPVoqaW3eEa0GE9vi+dVhqHPjU9Ujpamm
Y5JLomkvvfWNEEkMT2NNay/M8+tun+RV7jpC17dp3TPNtLblRD+Js3G0Dqaiv9QeYl77xufTXa0l
RO54LhBbvJuSJoeYPW2AeoW9OXbA4Io+r1xC/NFTPhvUsQs3uSP1MyRdduTwmCMf56UnRKTOSm64
6IJ2iOrhDzgaVEQtJRn6YSBgePnYJpMF9XJWfRjviAixQR70/4HMSMdEfz4ta8h/6T3E/OspVDfv
C48FEx2PZNknpK8up1/Q0PM2s4R1JTM69wBNDloTS6A17h0v/DOOwVJQGa7t3ekY8lE+1X9m7dK3
E3vN1h1kXJSL/13yWn2eG+/Jqbup37GHe/UOCf0wIQOXbfq6aQQnY+/6R8z8oG1BnixmVhGTPZKk
0FmKrBAwX+01CHfKeYyfoKfjtLel47bryWE/vPXdC75F3C40ODku0qeGaH9ONeK8zgcLH4wAc+Q9
JiwIHy+BcE6uDpNixQldbeKpP0UQ37GgLLXgVW579wgaR4aPLbxnhB5dcGODpn6uPb8pZfwGhG/k
s+XbRsljAafWsLW30GvESwT6wg4xdphVsRxjE8hRZ2dBq7pv/wcflZkedPbJzFySgq0HkDpsj/4X
i9SwIGt7pxkfst4UXn44Q5+ZE9gx0Wk6287flfxkjLH4hG8BY/W896jtVyl4dyq5aCXI48l8BXWE
FL0L+xufiYF0K3KuDiZYw1UNWzel7hR5lNReFN5KqRpkG8dBGnQ8kd66K1H1ZFEH/UsHTT8smJVu
EFysff56UsxZ3aQjB4w7xTPbShfEbTpI/p+N3UQMKUjIvG8zB+OBDVLhOYs1Jl4S169kz0Y1pqco
rZn70WYCQRNxatXJVHKc8iCbnax8lqNdqA8joqUWsH6blC3gGaRIiYGVnl9151tODy6f6f8aFyBE
DXxZN6ueehEkUjpvNOFq3LOLqkCYFmG6w+VT/CeY1xS8SVGQNX/gfc300KjDTgShy4kdH1V+OGWf
7umvpgBGICYpHm889ckpz2Yr+r2lmvNRgbfacFnzAQsZtuYoheKP0ZJadw3IX2MlOUG0sGaDR+At
/cefKF5AKH8WEJtFJiBTo/1U7pFg+ZlTNRfhsYIN3hpR8mh+5/ym0C+kJzV6nLmrFL5D48X4aWrK
py/+GspIJNhz2doDZtdqkr8b2YQyHkHeZOz5jSOTu9RoP4Bwt7g3/GgarFUKoOjoxct3P9uvLjkW
9R/8cOsJOriekoHYZsuR7McaV8NiirTX2K3ur8Z6fWTQT4ZDqf92zcAS+PW7xMctpNbs3pe6x2VA
jn+EJQnyhF6Ay1zuoEoDoGMk+NuNtE5LO8tkOBd2+JjgD50YPjW7eRBQlNHYkWKGxP/Q/LcJf02Z
o4OjQqg4IAFoIyGDIa31hFhKnHwZ6656uAoUv+XwItj+18sh1gfOFy7fZRcL5VJIbKK7cKpKq9tD
BHcEsKdT8J3gBEbeUs5EbEhhxvHqFqM4BC8eKOdi+FiMqI1sXWCn0JsPK1mDO/Y0y48qOwNTs+Rc
dSY+PLSmLjhDoNRAHe3oPwtSxWnFQVp4LTH6WoLLOLLUqiQ9ucqsWh4Hcb4yxbXWlkgXJuqw/4IN
7X2Xgn1cvhFPXmcg/ih6iWmnIrAGdcrsQcE9UgiWWxIYJO5Bg2BdwVEKDIuVpLT3901Z/1TnobfK
H5zzB9Dbd2PYxMs7RIpb3DqwGt1t7TaFCEM1evzogZNvpA58U8hHXwHVQH2bDAKfb5gVOl8Ocb0L
Em2Y2+CpYqFj7kpqUo4nykmaDXuOJVcwk4Wbd3+miAc0EZzw09vJ36+gFU8R8A6NAGL5eFVtFjPG
wXtD3VOcRsa4NjIpEfdOKFDvOtYmV9F+LIFTdj/cuxlYG37RXDVn0mKNG7HNXi4CLmJ1FgUeC1H2
aOQ3KiovGCCSO2N3H5rg8Ws3ricK6Q92/U/PwqlPk6lPHO/ROG5aJD3RFUWbyC3Bfiu4wG0KR1da
wBVFmKNTFvD+Lkiuptw0GMR0cPC4uwbxgyEPc44ATY6dftCPtRIv3W+GFiistJrSTcwozTpe0kb+
jbAS7wxExyz/nshp7iIwNWTSYEr2s4x69w1AqCBveY1LuWVaWAuAZzo2p2+Va8ggY0YwTuLF/IbK
b1kvCJJjZzR2KmQ66bk+OG0X/RL+mPvecaul70MNUtzX9OzCOvqfo3S778GzJ9PEAIRabSsKibr/
pLlWPOngcaVUtVD09eyMglOiJ2RaARCN721VY4/9CnKfOP/jGaxzZG7Etb1HVHlJNJcO25dTazVr
tfCaQL45IUR/7+RP6kv2pwzak2MPKBfLdMP/MCNhSVtIG5/UbG20BGbBhwMDeq69MZ2lwXgFMM9T
VS7xfzaHu8YYdgCbnRZFtT6mADBz4k5RzmugkGUPkyCOIvzwIR04aMMtIFbBZY3EzJFiwBL2l7rN
doJxp51BJ9C4CHzkCPVEpwtq2vKBgHO3zHPELrDrGqVsLlh6HHWMN7A1yEUn6bjKx9RbV3sPrIGE
7eM1C8i1vxZB7neeE9qL65XUnq1yS30fkmoA4EBOUzn5zz2XcQfAzhGAxPfhw/aMi1lLpo+SeHJU
Bor6Jsb16Lq99LvqIvfMhfKxAR3mgOq6qlpfrXG7EBDyi4QAgVXfBuLbe0WrnotFr74PUCsVeWNL
kmJca1FB3UiG4zBkjuSGR3I0CV/EhiIxLTfilZB/69FSxwHZ7Ycb8Z8FOaYKMpqvKi5GA7LZg/9K
uFyYbFZwX/79QCgpfvyEKEOBUcnwzu0Qg2a04blv3LPbp8JFpuCAt49V/guaXpbOKQyLThry1AD6
p40OUb71hJejrYFcnEaGpAwll6PdM1d4BKYFHOs85H1EN0ePVYJ+mLrhkQXcklV6tuiXdyRRBZcM
xaRozzVQnPiLQzfXvnI3KhRwsU1gjkDnNz8egYPdUN4UY7QYUU0ijx9baaU9Hszuc6m4tUqRzsgi
1RKjRrxZ0ej3rv680Nr0fwGDnCWeT1bws0Mk7jTKDi0TXwst+2RjBT67cTSE7f4byb79jLw6+5ov
IvZVYNVaV0hcbnXao4B0N2qJrk9Wu00/F8jrodFPgXutVhljOHJNOkvAd4RxgO2JmmBOGZowE3yz
Aelm0CrPKlL6NnqP3kXavUyLVsw5MPjoYy/ybOFV0OnFIYUOSD2tXtzCGeA6HyhzD7TQ9fQD5fmO
qZIg6E+VyN40L6CKdi4hoyahfX2vIYNkIuj+2/8K7IogoscN/5PM7WL8+08eJ0sr6GJQCE57nC+7
qmsbIZaxfMA5rSNlK7kDtyQ7fheoX98QPsIqIZgN3C3gDWxv2KDeWTANj2Z1dcMbKYYTBcsWZ7Ms
SEF27upK0UiirpcpvRuG5p3HzpEvcZwHM15epW3ISlNvmVDVpvbSXnltGj+hRODcT8hJdOGLOwnT
nVlAYUkUt9AP9aTyKY+Xj2NJDsPWwPidkNzGc5UGK1cPomLOWNnKP7HU0axVC/eKmO6ueUo0hG7a
cVKGHPtHGCY8JoQGUSIj381Bn1pS80xosAUsZ8eaT0QvwgCvZN7vDZwVQFME4ao541gSVTS7XOsP
5wWyIdkgaajcHRX89lWc9guOSS2G9TRhymncjE6SVXw35fRqdR5JA47sn8FsMPbPfdxmK/ZT2Wc+
dyhmPcxuSZ5kiIHSQu+TMA5nK6uScv5axXLyivsDEwKFxwwK0HpwXxYubjVgXVaUMjCW2vPLK1zb
LBZeKSA9zpE9i8YJBi8uvm2uKP6X7WXiahFYrC3LbK7BZnVeyW0y6tx4tK0/FFf7Y05MA9eWvb+z
i2gaOHjHWZ/o5iF3Nou9HDMGRgX1lVZ8cql3P9Z/+iPShxlZqnBOUB96XJnoXYptdgYbzK97pQBZ
Jl4CW/ReRVi7gsFGAWC7pq7wd01l86xlmJGXtBArQT/L12Q3b8eyHNhedko7hjTXTC6oR0NGGccg
kth1c5eugbsxbGyunjL7UlBmyj1BQMrcqdxABTsd7uHuzbYpb1UXMwrGyeZ7VkcMQy3XtEp1Ry2M
gBK9BO9XyWe32bDoNnJkYDkufTOeTo+Uv6Knztj+jyuLrM4BmMu9AjVfsX71TvvkYvMoZOWJSK0e
tH1ORdsrCDVYpZOWFxmeMxj23/u2Xkn9ohfNxaZ4cgrDIAabtsBz0uQ6sb2oClnuuJmswVFyvYUk
LK1xAF1sW57PAfeVSrMv5h89nSY4SzmUDB0V4m7n6jCmfJgeZ1dKKJXaaLqHs7GliPuWh23msU3g
cAqOd9fouj43/S1TxLUf9koHR9arEH7E1uCMDQsEZoxm1xr4qwymS4zpwVOHF2Br7x3GzoAxXG8F
3C3KXH/8xS8scOr3jqhkiYUN5kt/xSkndHxhBDgTeAIXT4huQWngN10cRU4foWCKZ5y8LVzkDCvU
JDeAFwlHaDR0+BSiI3wlKAQaIr1ERXvw1Oau0lcMjE1j4uQcB6HPmYy0ZfyOg0HInpGKd7ybNez0
ZOL0E38ZniDNkyNqjqJZVCSwNHws3roHZ743dIkGquCZ2GVYWmieSi9fBTGaRMeDG65dKeeDg+sK
n1kVRlNsVS7GBTwxcGrAVqBVZDvWeWDBhz0du//TKyfli8u775/IlfB/kLINdWYmOFe/TmKj0+vY
1/S/bZZR2PmjnpfzqUALkZy2M9uvG3I4eZlz02D68pXJ1asy87KwDiLQkkBjUX6Xm4aJdR/V3iUU
LzxjNDYOxIOknrcyEr/JjELSqMjc1HKo7wIQfSocumD6X2WPRtXQdYEJUkU8YaufupJDSKDVnINV
n9TX4OQp6abtIf2jeXszgso+kLrdnAAsPy3hkHtg2K7vCaoDJAMnDoCgbHGgMq5leGkjF266V+1F
uY1OOeXqRaGYaEQbAKexCp7hljKKpa6UUmFUof0Mjme+XzxcDX7iwff0sKDTrAT3fQV4/ijraVyH
S8KVk5xf5OVCVzgGGb84vRi3Zy9XD6PKLz4t0aGw60YNtttJpQU95hKkeO67Li+mMoIeq0g5YZLZ
c48Uh0J/jgHkZz1jw2gkKYyPdSianpDfIUHQwv0q9uGA7TETasxaJqsH2Q7BoGmjaAK3CJDmowKt
84DQYwxTFD8nXIesHF63n/LBqeCP1ASpBoe9VzAKZdxROCZKKk+9JhQGLgFVfHroPmJGq2zlA4qQ
sSYguWnJbiiwGs4vlkWjDQqdQkW9bIQHKY1AcldNyxJPa0l7a/nWYYh67np3ploAESDlN/LOacvV
XIVauCZ/whkmytsStmzoymoMft0CyKvt5K7xN3J2TrGB2NtbTxwlCJAQnuKL+/Rm7BDeOOSfHDjb
W7mivsUh5qqgESTsNXxWNtrpTOojSYeVjMLc478DGBtbc8U814qGVLeqE1z0h9gevF2wB6Pr/LcC
ITfPq3W6g52deSpdSvpDok7cXGjnCh0wWYyI+D+oItdJh8ePNlKC9occrooCkRWNXXQ8bOfJN1Hr
MD3YYjFulzy8eWsTyvtGOI7TIfzN9g0vbdyTPe5pB2grnJboTadzltMkDMlFZs9ZzH4JTP4wrl9C
mfyQ9VoqXfbuLUPTZC58fkXvNbtXkm5buVwSNeNtE34PSv0GHy9jK/V/WI642TCQBeUhtiPTW9hi
l1q7kwCfVMlp7OVBg7B8BgY0JV1mLSt0wN9ARCO+fIk4r+ewxgTggFJj1MbHb1a1dwXgYUSI+nSn
i3UDIdBS8bJD6/7KgMgInH/YmcStOmLoSafP/iXz3FT9xnnicgfYVrYL9ro7Oj4KZkxINQtRkehd
f7PG1EUx7IxaKWkkqsbvoeru2Dtg3GaPsFbWMvqgjROrZi+ntXDcAk/COiYDrqS+3oJMwZrN12Ot
xiAV2jtjGflLvtU0UWwvO6vf1ZXvwD40YqkD0kLV6bwnJ9AOiMTdx4eH7qrYpEM/o5HD6ZCZStK0
6SweP695202EBK8Tsn1IyD0ALIjOrME1w7lxqQKfA/bs/QXmxBmzGO0jdGJm1m85SCprOazyzQa1
pAtWd1PyMCzHgZEZ6yOvZeptWs9SZnYo+nMzpPZyT6ILf8PbSQGuJ3xtyhYNff2tDLeYaoQJqTdL
EpVWRX2lFknm2SfT1iTUmV3UegX5VMehkq0A1JNwposRC0c2sOJBRxYUCrcuI+YNlowSODyR7IaP
We/qweIhUfI6oIW+f+4capIj21eAZZE1jrE/VJ5TJsx1WwVF6J1/akjf8JCsZvXDBQKsjrNku/IO
NO6lLEcxl7aQOONRbH56NNSEvuHo7AUE/4kWqiaFxBrMZfoEUv+Y7NNah/IkThUILTlZkiqstfzt
gIR802cPL9uWGmeO17x7MnYitxAzxURr1GP/5ZXhG0UpsZje1MOB+P3b/yvS68zKVRYLjOJYaB2u
/pBBfFmXObahQaPAAR9IxszoMQrVLttQrxBXS5uw88k7/Q39mna9WrQATlUcgL/eaFdeCoqKW0L7
j8lAU8es4ZiM4g5gXZHAE3AYsyKNGRCfIkOosUjA9mXn4OMqYMvbV62wuKmen4lfQvp0pCNquiMT
nGHvzdKois3ySd9tejgmHeYI2+Ovn1lfDsaCW0Ik32gCmWtR4u3yHfqq853gXcYW9hJMSbxBlc+d
PF+rBl7a8HdBz6kgX4louIuYqE/iwg2ir5xGlVxywDDU2rwXPvG+RvZUPzsEquuASQDGscFYGDQH
8SldAQVv6QfATiRuMJA0GZAvUcpj7yxnBIB8IxPQYOdL2wzdSOnFWYoCKBnBbOJi5N2FNTe0VfDO
5rbO35Lntt7hG3J6hIVlvkhomm7uMx0m80IXy6ubChDb1704lpY7Oki6aNHX1iGokaXQkb3mXKAI
icxJvNuXN4kfpzzSv24lTfjMlNuXIdp5y4mWa4adk2yx1KE5OR+h4Pc4aHA3G6M1g2B6x1wPxKQ9
lztcIhkE5WJ5K84XwndRi/255YnjKtANA74odxaBqZag6sfxdIdOLQnzRbFtOXxXY+10FA9gJ7g4
LPnF5U1kKiI92B6+z7feMqPn7tP9wmiKeRQ4Iz4ovDnwgpGaTNtXt5cvzLcLwZEojs5sLG2Oz8b6
icsBfqeB+bN1CBtxO7JaYe+FC3sSWVlBZZP60LsVSdHG+oPoBxwJicG4cuJcXkYnN8VMyDMvSetW
dK2i8R0Hk1Eo4FH4BF6ALylM6ujGCk+m5Tlqs2tqU8uX+zSR4gIwGjAROqgV66Avelef+VMS0zTV
bQjUUN/Rj3HXtKRKFAz3xA16wPj31L0afJr2lYhkqoHAZN7Or4bMZHLRsgkNA7g6sKPngzP3OvZa
z92jccsbbv2cq/5SelbUcr3XGFZFHIcwQe/suxWRpH3gM8Ubb9hmuheIALWnUgoSZogPfzjG6/x7
ijtQ7e9A+gOC6DikcSZ31srTZA9QlM/EbwmfucTAwTPurZeiXjROdxNVP2NSWD7jBDdxvd7XBHW/
d3tPBdqhgAD9fgat6n78B44uIvLPjJOSMPW7nOBOSlxHxYtyXcwM8RFisCDJXmZDmHrVzb/ByUtW
+FM879U52yxUL1uy6lVOkfzpDXjBDbHVGIV35K7hebBxDpYGwHTmV5RsllzDjxxg3S8JYR3aQEXf
+ka+yOVxCG7TA+1kjHaREEVl6ifMH4hbXPwHoefIwICzzpTklter3mUIVrokAHO1eoblgxRdgRp/
n6WtXmKiOfYqOsRYyi2sEdS2lDOyeJ6IG1zjFj/v1TkJBMNHK14ditFhl519l17kFthd39uB/LKr
2EwDfvXf2hVthMAD1m1G5rVLm+6Pf/tFZvkTWXRIureSlzJBpBJubtmpuy8NHmq9LM9wN9PjhlAh
ZNGFGn9w1WKK++La/2pGgoXSZ3cR27F8pP7RH3CEO3NZpGRNoUQIsSzFBkVieAhAfaUCmxoC16f4
y864Naik5sNfLEF/O/YKucvsrSL4/6BW+bt7NCKim6iJd1KY+hfH4DWfz5ZdyUh+UrAurTrhJBRT
zZCBVvrCcYOFoB4pYOr2Id0YUZJzq3HaHxo7x2rtbF4qXMQafYYHcijxGx5ujNfBTdYaNrVUYYBu
CIlxt4CwSH19nOJGs9EpY9dL9qmRVf1tPfUzoi+UIf/qnZL5fEavVioW3buaaZyhD9rS5sBDUHEI
HiF6Qa0xFj9Y9duisx9QvvkWLCu3UNTBxVvwVWbyZOom95/A5Jkgwz75fcDnWagPrR22fFYJ2kvy
0xdayOpXlw4uPYyqsSub3x11yi0R9mZtdo87y58XkYxBQHtmTtHzsZg/rjEZcfh+lmXf6LmK2L6u
yjmwjQkSBRfHbP5ZP7PK3QZYIKl3Sx9W3IIRbxOPRxh9EZDYTDnvNwrpWb2cyo/shM1B7BUOycdy
lt/egasoy46dc4ZR/5Mex4rfAhQuXSftbuarc17K8r6jhMhY6dfdqn91xZ6v8FssHoF3a7cL8tVg
9BmoqnLRumcDxE7mS5gzwIOdIJfPTc5+Zp7EfT3Kg5L8AL+Gcb/YHWHASKQ09/wdH6d/sVc1tTYT
1J2dQ8/xhdIzbqYvrFoGTnlE/NSoVwHbUYWTFIBuLxBbUqXoSu1ywRR8hanuOMhKhfqrGZHyOzlv
uUBrNB9OIE2n7B0p8XrJ3yUEN37O8RPVg7cGu8ZLxxZKg0b7Hk0QC5LcUZZszV0n5lEwNUDmTvTt
DWttjmf63SrGstQgaPKV+gkxKkmKxUfse1mMQ9moOJj/vC8rl4HnAOJaNWkz4Es6+iEbpncsoup0
bcJ1en8F5nYJ044/6lZjOJ2TzXeundaIGqkbOWG63gHZvgHRbiRZFfruC1z3FqMqHgimBW3Apt12
obVm7zoIprTQFfbmb/ZEqkbHWA+Q0gydoC0kAzpk4+0H3wJ8vjM+Jahelk7le8K9pcl3ky0s0Vlf
5dEmEIJjfKt65XnS03NUf+mdZUuu8CZuHBpJfoklgQY7tv1j1NWOKLWIOrjlINH3PsbKVxcUUra1
CYFmfQreooG7QZW6JDxtAJFNX0O/n+ZrZk4xFgoG6lCZQo+K8wXlmDz9IjonNOl+CrGdmS6vrTUF
S1f0lNofm969a17728lFWDd+kDWCtcVxj4B0TLV9Y6UTRpDdg72PDiUYTtXifW6WE/f8LXiz5rRv
GISo+PXs9Olgb+6E19Wlq1uvEcIvBqYShgjf9JxgYGF05U1IlZATGA/OAa8LBpDNceXskBhT65Wv
uay+EW8woeppfs/aa5VoOkmtGHg92ZrfuljsKxyxkISVTVbmQUwKHO//unQHxzB6La+3LnNytWLQ
KwecodJQMA7EVYzzhoLLjlR5rY0UrPme/mrPJPyk3LDZIszOa1eiR9CfdZZluu6MCy//EMCIEd87
hczSRCoZ3cKcchc1cPlL0w8258TPaZtCN3Vz63bkpgtu0iDHFX/KDS7BLcnLaj9EAg+xbe69rzyu
x3BYE3XiFZsBNJbFaPgbkp+n4Zc6hkVVPi8QFycYdKPfRn9J5ISYLOPfBB0X5CwErtWTPNfF7tTc
wqvGEwujLIbgioc9eUsK2jCKbC8IJ3ldQtiiQiw1DRmcCCdoPrQKKW1wpdkGcKDDksIOAoOA6wBm
tbAD3hL9IxX97YwNtdns4sU7JT9HPauhPQcO/S+lLM2oM2v0v9hoTAWa2R23RfvpKkz13U0uytxH
h43PzG8Zz2XFOu1HCckURCLnPBdRB3MdVXK1LmjVTpxXxfT6oSBpzWVmxuoMFQphpfCRX07TxgOl
iSeQNDx+JcPNKd6TlzjvHYJKFEjDYVz0D9Zxa0O6z411aXBxwmfGJcvAZJsryW/4GmMfhckve7rp
MtICZvvAv+5TlodOe2q5oQklkRVQ1ab6ozcuYGQGYY8KijLnqRh/Qv2T/sqPXbRd3raKsSzNTZ83
t3k1AA/bmjSJc6hAW1lCc1ZhPB3T5yBbt+Qhb/lLbXlZ7jl1joJmjgpDEnJFHVPnnMuEyZvQJzbB
gafMk8hqx06PcBOGkMVD4cNPudoYq2qKM2xO4WuiYrNIVhLzJZDpYo9mHGekBU02M48iyKBsDdMs
yZAlbtfkpIF4ypH81c+gSw5KxI8YroQGrL6fXXuD/yPekOgujaRV2n6ktR8jDaKw4lQEHOwrlLU9
9jySVcPDbmYjLqdz5DdRdw7t3oFAezFtsBjF4Zj8zCtTHf0lW9DTGnqu97MObtnhANSR5F54VSXg
2MfwdrpiF96vTEQK8OOkhzpTyE6+biLix55kY//YwdkDsPF5HBC6lC1y+xnwM+DdN+5N8JyJomac
6BIN/qGxHVqbwNz6QETo0G4SzNwbSWIjJEM8LYFEOHKqbIpTwxGaEfQZDsAOHjXzE5lQCJIXnO/K
7FH2rAGznbMZZx6DesKD0fZW0MyINq+s8dK0GXxAV55PSYT0eyLMjIVcfMZsGBDm7DGEDKhw3ZL2
gMesPb040DVvAdKRo4l1rkKbjQhZUEXCiB21c5U5Jo2ICwGhtIwy+qAjrku1zH1R8l1dum6MID2H
MbFrooZFqghsJzzHYHhyHMUuynEnz2paECf/BXJ4z1Vw6itQlM5HoYUs6dQg9cz/qBCf4n9zNV0q
wkl6nUGeiO0atJNLTrO9mwfPu8zimZNiMRIii7n1jN/P4/RS5mEVTAu2V9TATm0OWmxU9nuaWoFQ
J9Ee+FFjVUAVyz1NgDcgjEdFEAP8XBaW4uxK+aI4NiF9LmS7jEpVDXD3vzitOdKKdZTeKNMJWvnQ
lUCQFXMxtj5AlKKtzUVmV6ijj5a3mxIwlvT9GJmkfoGPNGRtxiP5LJfkEJqf5CCZDGlpplHqz++6
bSvPuO0qumj2pIFiPn27J6dnv4RMiSb8RvcA6LY1/V2br58zabV7GGaEYmQKw8LBSyBBsGHMwe8n
gvtZl5YBSwIErtXt95KgAtpTs+IEG/hKw5MqMP+GomNg0En8HUr92wspKYhuKBRk8TIh+3+BSa82
dVdwS72OrjzDg12Zt0zU7yfEif4XNLTxFkHy3UDLqlbPVp5ezXMsfI1CsL4VxcmdT3rFfejUYr/T
TqXzJ20ohJ2Ay6/ZKPd/eHJ8eAkKArZiQIAjzvZOxxYhwvwrU1TjY+G+4/8LdsudohmohIiyebto
lgMNBhE54yiRicBoVQrAGfA1mrInFFq3cUMIt69mGTkYGDm+BXNuldrEdkwuoxuba5jE8lGJ2HU0
10qQlp3qp/54kg/Vz+sJrQZdB//+4FSKNQefVs3Ixbgev9/Qfp+bupbExXUOIH6TG7I7xipyMUbO
RNl4yvcsJQL+4KSNE3Fx9DxgZw43A5ZnNstsWmMCz0iqyFqCA9t8Vwk4C76vYJpRyRIAxYi5l1+2
TPGPTj1lXn/H0D77fWIoprqTAh5RjXGSHVaaPpx97dbiweEAEO6zRAstztJV5Bz96pjLJ9tsPwu+
5Om8zAVy7RLr2N9CuLIBmeAcOF2VVwf+Rpzn8817+xz2iPHKPjdaSZB0a0TJvWbCXgnv0YH0tklu
24P17Ov2gyvsE60c2pzmpM+5N8E8Z+3W3EAO7LTuVmgVJwmQy39Eg5A44hMef/TE5aTwKGasAWi+
jRHuHDWId1YG+K9Y/WRfy/Ypf4QW7bGUDtdTDfiZwnYaAPm7vW+deb+CJpJlYtkyYmmkAyJfPHVX
ELv+7w21eYobwwgYog+uqbTlaW73dQ0Ex7XToUzglB4AuQxxXZ4QpmvyxdOP8QEYv//0V5ko6rsP
m+JpXhhVFEuwgpQC+WXXGPshKGjYAwYIcchSXQxOp2uk/jCtqF/UbOS7EgCAZu/o9yR6+p8Z9ghr
mW7UcQHYHJ+FinzsoGUTzHdeKPdgAiS1VFZbrHMHL0Ltt+qwzDTvJTH5X+xEBNAwU1IYs1VCZzFc
6px76ExFZ/BgoBR4gO80L2RdagFpU6H+vqCGipEPT2MXoTwTRbRgRaLzERDCtYLuXvr/p1y9gKZg
XHuzbYrMr2iEzz8kEx2KVZFT5nhQOgDLF6egCsMl7yk7+kf9gZLryQ/J5TVnQuiu6rgf08scweOk
al9LTlYUK3sjRcT0EjRZpPK2yfcoQK6HofYxXBHo/TbOul55pWIg2YT6AGNaTLh4hJlP0j6Ti9kv
W2eQfbBLCxct2GF5i9dpcjvF98ZldwajJnRfjz3XNvtu6roWNH5/9x07xdNB4mWiuoMEW4CZ7E0a
DWq+ztOQiCLDh6FCODheFg4szqDazOwvHJ9m7ucA/uY0vg1vlLHokbzu9WUjEn3XqJRbyu4aoKa4
I7/ZioVAGv9m3wiAiP1wa2InUSgdE9JJqFEm8cusWGy8jEqAGLiPHeU1L2z7QplbFo4dt4XVNeYw
Z7sW/vjrf4cZ6E5ENJVKZ42qJ7k8W9h8WJZAfmhT3hAYnCqrkv/WZo/B+RaO1T0eAhvpmdMYXOIg
vStEBuuUgwliXEzM19QOviDIJZJoBQmt02W37Sd+JPwl0MaHEawMlH+kB8V5WFR1JCvhElFmJr3y
XQgxgxULpdPEsK84rdFHv47mz1A2MLYXbo97bq9MowToKuC43RSc+HbgYneZmV7vHUUVOUBuur6p
7YWqfZNZjPZFy3rks6OkPNHJbSRZn34EBc8vesRLYWaCASQpTm2WKiXvvM10jo3KLQr7bKgrxKtl
F0vnya1tqY4/CU5VeZG2wC2KOgOZ9CmgfEZvBw1Rz92ZCJ9ziCHjpVzwChtqwAYp2h6DiGuvP8RG
L6BFYhJxYVd49bgzc0vpJgwOP+Qgw207T0pBlWJD5ISFujc/XsTwyJdrEvqs2sWmxDw56m7/gTyH
5kwLtxE8nSS6S8nibCtrsCYlBaIOYl2EYEOnHVyyK5X4RccAvNeu6HEZS0dPnIY6f+L3kr7WG2L0
xJ/EJehUG7mOy1pPiTY+wCbumLoQVd47Zha9aKkw3nGfAXlfwAo+zRYPIK00Y3WGjrLOsHtMUZtO
zZnTQ3LI3pWiwIFHwBhVfeLoWtzpVf9Al/Yiorjn1KYossFj+KUVQJnin8By16gcx1B67G3GoNlv
XWqLw55hmoa2hwv0hVxiJ4mmfcBgnba9vjE+txUPBWuYoJ6VBKLY/Gr650fgTgfot8T4JMSOyphm
51eBqfpIiVr7jWmt2Qxy+J7SklhRyqLqyAiInus4swHZZruKVPG/irXR+cubFzRqmzwDcey+b5Ph
+8iTMgjbjNBXng7z9e78NKjhOBZbgHM42QTZrAP90Ql4UInEOxU9Ga8w0W6DvL9LQLE4BAXh5mT5
lFouJutAcaRfqBMVUB4nXMTyyh1IPJZThH/PCDbQOmPNNasQHw4Zj5GYqL7JDQvp5gj6hbXbiaOt
xwvBs3Inzc/1QggUpSgo+ESFwAl0rsfn49eecncxdFhLUkoXwlvWWLVHjh0SSSRtf4WHHmc7+faL
HwBh9gHNEnl96KivtoJTfI30abl9Xfg0CATLZj3dFayhk5EAxQK3ew1SoPIAPhdIDRvLBwaXwR3o
OW+oNwZGPX9VfZSBgduPpGOvd0ZOBYzyRTsUab+y4/M2mCRSPqvI3zIIP8GHrSyjN0ZFGdFGlvDK
7r/mBP42l8hxgwOTOt7OXQOafzwiUGNr2H4DjQkixq3LO05YKqG5evRoWbaogoyVWfesrA025mSC
wpHgD82hO7GLHVHl0s4vaI3ei4I/l4irsLoI+Wni/KPcTJNLN2GR85X6ab1NDEL+LFVkOlFcygNa
eKUQbN2CGfyz9wA+EDmKQ4BLen59uP/XqLxQFPp3ecMEu6qoD6TjoPoiM/d23oPCYLHwq58eF8v/
5MrNhJmzDoMzcW7VrfjK4lzZMpy0TkPO+hJN2rnDFtwv2CCmjo2w3bKMCvS3gjlf24yug5F1Gp0O
VcHaelI0qQxtecySGs0zu2MorI02QU4pPCGtzVJdiFgP23ifDEZesyzzHvYDC1gAV8zqi+jneKuC
6Iy+diTy2yvGbSP9sM+NR40ugHReTGiwrKNBWo3JPAgh2Rj6RNJZ0CDWHV+dd+R5tVcbGG5NuWM2
T5/mlHWW6RMWKqWu9jxu3PpgJ+CPnx6v1xOae5+Gu6aKKg6aWUdgWOftrTwBc92NAj1v8sVn7Kke
L+bb1FCTpVpV2LJci8prS/0VTM1iYwZxn98KuJLtGZhK0nu7y/bIWm/cY+Y4Nr4W3S8GU2G1O2JW
GSSigxzN61GvTuCABZVZrpskxchG4/xf5kZh+Ra0O9aIgWH3Ru81k9kvnlyv2pteabiSdsEWIpFu
C2XOEpOSRx4+NQfK9e9AzYLQaKgKhjwCMt4tEvEVaFzvTjj7atzMuF8XeFnbDHj6oaOYn/jJtLgM
ON1KClmNKI+1c+LctuOBJg6ToGrcUwY7kcz+0qbahOGCMruYD7Ek4azHAV8zYQMy7pXdHPPQCycp
MDyMz752+iJS48DKTZRA8pNnycZLE0dbFGFdjmSJsJc78wC6MwxhG7L50Hm6ALX0IJToJ4fONBiz
1bixEIMmBLqnuH2ks/sZbxUu/FlDhj0Z1Nwn1FQtyyY4yUr/ucnHPrW4CC2icS7tcHhEznsIqkVt
ewPZH0dFkCAhY8P9lcl0Rj1yW65yQuFATSrHSIKg77sJXMMIDTU95wGHNJqfKkZrwP2k61GHG7Jf
k94M5T031QFt3Yf012mPln1jG4rw7jIvQr77+tUPfKbCV+oJ+hUriXBmNXivJ5JwjrMt9hfG7aZZ
mIyKr3PLXsjXeBR5Zw2+s8BjxbCyqEUINwAl0etHlxGZlywxon3gmIEHV/NTZaaXwxgp0D7NUfMf
ZZHGH7DqQOx632HOyJaSmwZc6moX6hXfjJ+lowTxOsuw+y/LsnQUEm2c1pnQkCVuKT34XUtQHmKN
wjLDN85owNOT8eEYCDrOmIZZgLSKoBIN3rDbSQnXS38xl5GKaREIptT7pPoavULttk9BvpGuU+fz
aOaC0HU0UZLx4qY7DrLfTPF672WZbG/l+1FRXsAroxosUKN76Qv3Wg2ONwABGYrWAs2cFAKgdoAU
oXcUwSvwY8RXsYYfrvYkCDqmJwAnj7wVhRwFFE5QDi1q/M96iMO2/FF/bpnWoueVtDlILPeZT53G
PNJpKqAjBAXu3uPEuQpya+nmi80ZHA/ycClamfo7MKHBkvzzF0PfPx0sPkysMWjpqblG1IIEUzyt
iaNd1xIBCVUJhh7M1QAdZ7AUKfv+Y6IeS/LYnPlz9OGkZjilNCl7obxAxQCIMqiczRMryO8krWC+
06GoFROTC+j3UN5wH26mQ9DEY6ZJMd3jsbv+Ruzn5/6KyFhFRoOzvp7vSdUDSBw+0lZqazAtl6Un
hKYB4LgPEMQzSNIzUtMf5yqf6KIWTp1718RqmcP1zWAdI0DlAtatHDW5rfsCozIDf0po4cfayrY/
d83k5LHqNcpxPORmTHGfAOsz64Ycb9xSW6oyqJhGxX1rJ/DLcWgokvNJFTHwJlTlHrR0yrsDNGWW
hAPUCZ6szVgqR4YHB0uVEZgA5Wd7S7amoEHJP2LLH9Mp2xphh9sxOb8ql2aQNIvOQwOf/84LmJJ+
Pt04DXKLjL4HcMGE287qRa0G8s4yMijQ/fpXWOosctIuXQWKxU7Q1oB3m7uyiiydbNAn6gVSsv7d
zYWGIn3U5bXOdB/R/0DZuZzZZTQSlbEPO0J9hhnboaxavV5uJbh6+9B2w7kyVYncDy1KRwPMKhfa
GSOu4p7privqqu5ToT4GSvPX+A960eRyL7rmQCzxel8/sMl+oUQGUZLvJFk3Cm/nk8Do9sDN46TL
xaulXnz0TaJgENGuWwIlgb1VrZ76LJQRKqU8X4RDhDhFR8Lw0NrGJ4QtHOC1J/agdFUoDi0GPr9T
RhwPJ8SFeNl6iU1rnoLfHHXdc1KEnCr7djJXgqFEN34z/y5bum2QoYli7c0D73oZgsUyu1lRVy4U
lB8iHBCaX80uEGbHc32aXmTzXeYcDIPY4RZYrsGFVcSlhgrBBpnYFn80+GHHQkT3FXZ+ALNQJVAj
1Uy7q3c1BzYn1Ef+J19DwBazn01bwk3evV8EMChUa6dJk5+U0ltlg79t+zWwHj/1fXknzBSn2mlN
LSenn5yy5+4RLg0ebq2EcfJzbcvMooN3y3lQxqJSFqMdGO5fL2AnM94HnazX895TzZpMqIBWSP81
sQibgHCOYBzFQj5YFXJMBT7BijS3YSTMnpXX4Uv5PHWL8a8aECNyOCgZplXZv6hlTj6LfNrcklph
g5UweXUOiEcQWAUI4eJ5B3MOtWnN1kt9yEinNy4qJcSI2iSWFOMsctssVZ35Ng88UKYzKhrcqDIf
W9dowVECLi4gHMCEL0DTLKhO6wWflqAGC8fv7WtQiEUnu9bxBrvJiwmxxOmIDq43hLiYyVY5qBlU
DI64ACTJp4NQOEGZPnzenQ5s+WkDtwKtwlH1OV6drVgQHuOn7sYJPvkuz8z0CejBUBTqte5PokXb
DGYaZxKtAsHacCE+N6++MJP3Hl7MCgabx/FMoenrBBLcWEZZoxTLTJJ6780CijVrVK94YL2h3/FT
GQWBqsxeTGXz9Cdl/UZaRZF8CylqimEEhQcXySsQv9etITNS8gRw8t/5MvCr5ajGGGnIzrdSaCK2
RtTS/KQTmon00YGb5dQMiofyvjvWOPhv2qs3R+qfOIh/7NlOczGcBrBXrZX/MADdw4vGvXEDvYS7
5yE+yVv4PUCnmBYR1hKHMKwmxy3QWiBIvLryVQFD/USTkfsWKH0ZPxa2/iKeSGelCM+p7HX5L8/p
C7Q+8TmSoIlhDELUrnhaeZT9ObnZpBP980KsE8DOyd1DocGep6B5kI9MVueAL34n36GjUAvcL2OV
s3nktBKvens+ApqXD6tmg1pMFnTT1qY1QGoHbrjKkpf1YJW84/6WpjZKHHknp4FIGQclq/LvWstg
qyK02XXOMBDmLewzvU18gTGMDGpUuUa0L76AgOK0a+NKeNgF8/e0eJ6kte+n2qoQFn5DCGgvOGlO
6Igs0vHpVYh9Ab2GecDHz4ILb6+k1kLvHlHdTyr2lQUWv219oCn0967ho8Wh7iZV6ebGgMQoo7iA
f82TpvxOpOcw0xjfadIOfP+ZmFUYFEu9063TWjZlkwNriROvOPNTRvg6lRASMPe7nuUDMr7D3gGi
pDHgiwI6qjSGSB0z1Hknlt3C3B74I40wdBty2LgIFBqTGScO6COAMppgyfnEK167hhJpeZqk6Vyd
FHsFdzIWqqsz9We3eCzt+O1t0mMrLyQG+w+qa5wAfdg5CK2qNUEBnhCbKXAcWdA7wvnzYrdMj5rM
n+a6lBgudhBCgAh2k4rqkJHcr2B6o3U3Cp9LyynBNDPc7qmC6zz9IFbqGg/LfbpPVynIjuGg59Ts
z1HOONq0qtCyImxV0Eh+TIcL/SLaDdIFlSQROQ4hV7TxHkAoGT6MaLwu8y6agOrfHjWSw8iLAInj
5L7/8GdHEv4WI0vKyoIRbheKTT7zFpNaLSkEGQcHuLUp8OgulSBsJh5fG3PZ8DLyLgffGNk/jbGD
Np452p+WYqi5F8gclaXd8EkTQyhZ4KhBiaGCNif6OMaP6b+j0gd0pnljmxt//VphJ/Mv4MCL9Pge
mbMrgRGQi1ID9aGQvDPAVsu/9KcUnpj+9JrX0RRuqp6+kxBeKTSwl9md88+nKm+QkI2I7dgrtXCx
elU5gZzurTjOX6UDqM6O40s1K2ycTUGlnvNznwRQDqgHacy55OjgH6becIHAe2/2QCxZ81PBUSaS
CGe0oTLwTJHKLIy5y7V4y3tr8tJxP9vXHKjaZMWK2Wx+6lTWJC/z9JlJZ6r2WTKeXGg8e6XYzsPs
nuFmypzOgexrduSRVpJzBynh6qSxxWU77hAd7WexJTqDttuk+DiOJbCQAvNmIzS0/gCnrhCO/jVO
SFvqMgttLMbGKEhok1gmk4+N/BYzT/mQJbHugk3wRPjJIEPDoNW5yT078dYzQdcR02SzheKSSTcI
d4TXQzkXC/Pb7eWYYAISjC7HmbL/PHIvarxiE3hJCjQLCLVEYRib27PJYRtFCVqTlzEiKY+Mbfgo
VkrHUUgWj/DnAc5H2+/RJTysD9OBAdageOcp6gDc7O/5P7QSHOE+UmGt9clIkwGb+GOXi53XiwXr
WiN5qSyulyVHheIB7gPPTO+YTsCCVLvqYn9sngVkMg0K96AcMkbC1KrQ9xxC0csyTEcXo7eZ3Gem
yiZt4XxR2QwWuXLXWCsyuRYYrLquPVG9FK1D2N/r2+33cAYZw/HqLosAG7J9j0mcUz/oRWrsInuX
NAgD0p143ciN3JUiM/FfaswY2XEaBsmOcssxJnPDHsxfQ8aFnfknPR6Hoig48grgX9Q+Kx+di7J+
j8gc4MBw9efJ9ESToPTAqLr86j0IOB2QSvwZlFHy1eEzBBxXxc6nIQ0xHmNakX1wsteL+Q0Ndm4N
EByzTWHEmj471rlcNe/81jInBo9Ekrgb9z3Qu4hQvJUJH/ClK5nyccRzk9H2UDbaEE9EVQcWenJB
qKm1l4LvAEvnI2/6zjybNLUa4/p2TY3ZxxfP3hiId7rNfh9nYOJCp8ggdsxg7GmsIldFKVMg6mx5
YbOT7vc7F7TgmUxM1a7eDwieegAPt8T0GvJUE80rDW2+F+w4RJHrqy1S1w+8MNs23VBdrMVBiso+
lufmR6SM58/hB7eVU5Tdu22fjcQMXYEr8XUBNT86qlefLJASbBCmZO2LBYwlg78q/0IjW2GkvTVe
LQP7/Cswg4/SqWA29sfn0o+CxKObjYVTWt9Yq9oy+ZWAZhMh9LU0QwDPFPp0yH9j0AY2L+w4D9Mu
PwiyHfznS5/eEt4iUj9iolhIcXo8ynqiCWrNo6wtX/ZMvEr1b5NLM5Q8tSoeOMlVGpOIjkF7ltCf
hFWnC7unf958e3U9sped57OWa8kbfRrble7D2hsSVhwTo9Bs66qfKwjei0CTvIDPGBwJSoQhW83C
0I3MESfOhVf3PG5C5vMIYWT/54RxUNnapobYh02E1SkuOapnLqfaa2LW0IfWwOFV0SjaNIXK2vQ7
kYCVWSMds9VP+3gS1rd2KUAX13vYGBZ4IQxj8j40uY2fJNdZjNyNo5sBOr3etEzNAoWPZ6LijHCE
LkD0/5Aa80NfZRaUi/6FAMsdb+L2/fdlqAgNaIucUEw6V7gr5o/QIkzJhxi/T6Lel6QCVOg13LTD
IJEszngfT29oRtTsoPAEy10Zfq2XAUjyxWY5I0JTq/b8BZM4y3K7KrfPblmk5ySB1kLUrPx5jOok
9P60Hem2cYZn1DGwXUbwB++a5AlMrGQZ7r7UAmEMgH0zWhnY6zhBgZPybekque/wNVfHau2InEtm
+7P1oT75xaRv1+fB+8rsm8Qv1LkoB0gB6iJRBii8dnnjPcJEhn+vIPl3dhKqjx8SaEsw9xX8gT0n
KNk7pnrhPnVtGv8NQnHLK9EXSl+ztrBnhUlKn7+ZQebN7lPqfBM8Q2tRGezRuYzI2CSWfLhSAXjr
mMoQTapWs4Y05J1qwxdvZHPGbmL5e1fSNtco3XiB9iqNzzoVoU/umdoFFWljm6BVvwBfBsM4un28
cVAB3naJlJnMwl3upBvCneb7nJGZeTkqh0kjvGliHB5SijDn6abrzIX5s9o1T7z1oXGmMKVlScvC
BSQOtCtIELGaY/Vs+gPo0Dm2EFQQPppj6eYHoxu5h2zt0EJ6G4y9K0gxcj9G358pP6w5MvFnCFes
U8QQ7iTjmjOByY5lYJRmEdvgHmP61EKbokLwv4+mv6at4CC7ipjhpxqnIMD2FcZo/yGKJY5zoziG
Lc1hFk8VIb9da6MuW6pclUCTNRW3dXIDLepwoZVMQToT9SiCFO45c7CKKmaI0+F7w+CPRHBbZZni
jYcDIVlhuAGXZb4iZVYlOukukGYaGL8O58PZp6j9KePJrJ587pb3YdJVJ1H7vSnOC/7xZATl+kED
vGTVsMvfKxJLh3EMY2Ngyqu6njKydAYiq3+JH+zSz7mQhI7yloU+D2gi9FcelFhA5R7Z3G18q94b
OQOaVLWImy4twgWQCv0dhyKyTgYSc9ek0INxZQ9zgmE5V5ad3I0sj4joZwaU5i0xdpJlnden9Zho
42Zcd/96guwwz7t6QsXaGyqb0pgJX7tsciXa9uwIdpSgA9TGnz7F8R6C13BznOCLI7PffK5/IkXY
H0AMDth/HJzCQ4CVUlyVMr5aZ1ZFUPVoP133Lo2gLHiNDMmOts9G4f2CX0j/mCuB/Z2ohZ5qJQaW
2iFYkbBEtMZZ+QdwHLcD/C5futRip4dhtdYKiozQSx0iES7R1/e+6VoJNl/IN4HiKguArzhxE32e
ijvWygaAu3t2hjC7MrhP9oDIZcpbXrEBXuA7MMu63iJeLPTkPco5dmibWUaVl7ppSY9Eechpje10
1GOsYx3jHNwosDxyVc813GuZAqvifbu644iktZHlTF2M9lODL7soV9+gMCFAV172q6qk8P607ZOj
zUZz8znloxHOoTkz2NsXFNIesRSv7atzbPcPjiy3JUtDKIauFb9uL0oj7SctV9q5dEuLocgawmRt
N5lDNjgd7XQubfFZzVYfexrb06Q3KVo+kNH4emkF14rUJBdFzf6r0TIeflQ2hJ3GEJOPMx6D/QNu
VAuvUrdt4k0WBATqANelpVrujtnn/4R8YU87VOhyoMRbQLkGDCTGh0WxleyUhsCB8abfswgZ5fUu
HoVIxH9z/xP90irPlK33Zyx2tjL1hpekvaeh1YtbnweB9alaoP7vQFdI+iq1XBfP+oilPFyENEab
pVOaW5askoXIjslmgE+7G4u24tSDt+c7DTc30uLxYHdsVhUVge40211r3RTXfSI52dDPOskqbgFW
yxVACbgP0fpghxnn1cHcZblm0IQhBan+gknZNgkkCyhtiPgZJ2YyJSvCQjJvThACDVLAqBrZ0hvr
knh+fwJEaP/PjZ9U5tV0S7bxaHqmqo/Yfn0baFE+td8/5ZAEkaVxYDuUWjw+vGxMEp1/1iGgYlni
KdZtcn4FAHEgvh7Rau5L6ypWUu36ngA/irlXnKF+bIFehxAaNlwOWfATyxxuhXoUgCck+kJvHfkU
JtdyDTCmiwdpcSrsF9wVsp51T5y07s3JvAHvL6q2C2Tmn/y5/0V4UylH3XPhcAGwqIno24N4+58C
Y7v0D0iDYvqTORV7TIO+LsNaTPVmW68QOR9F/h4UOrKsIrrpQ2ykYfEY5U7jRl2i3EvvWVeYrTXs
JJ299YYXUKyAatTqf1frfFnoksBHqq48TpOF0HMuJbEq9T78LiAO3oLbneC/owB6lmjVoFj1tTx6
DWRE+mTPdTdX34JMiLUmiBW9eSorvGhmeVGxKajEYHeU0eo2eUPxrrd/TKHP8MeEBd79bA2XB8lU
Eaaw6FBIcrlUjBXa3Av9P9VpzKJoQbuLqA3B2Cx7+y6UMcEQSOJPMvwi4Lpr6J7hw5GUEKK/nB24
kFt0FwntWEm/fQvz5m6GAOafNqLtsbp6TBs8awwOTw+T+FqfmAnwLqnW9bbeuzT80Cp9y0km43Yi
AN8Z8DukIQnSaINBG3b9vE6pvpoPLxdG4VArg4QWfJTEessjaUx/r9gdTP5GY7Jyj93tjb5pSEa8
0VsUNUO0OTGILVn6PTRFgcsEd1854dZO6blkLIdn/XOrVhtlqsmssgrlpXqFfYImtxuDe3kACb/8
x4VgNwRjY/ULKg05NQKEQL9ng1viFsZnSQ20secqK4XmPGlT/4ym9oUEFFAI0xsfqSvkmBziJD2I
aVAokbaygFT0fJ+WdA5maxXxlxxFNin+20RASNCSm6LSQYz6V6S1FtcT6JBEbRo6exvQ7a+IFLGK
frCZSAMB4GxnmfSzUBephJX/BgZpWE9tBv86MzJdAjDl1KmTGvnaXNcE5Cjv8NSvv+lQH1CuEi7q
Qn77K4of81YZ5R/NpnouWNdILScNUgdDV/MBSrE8ydxXfpC0BzFgDz+FdHK+MeWkXiRxCXgfsWe0
Q6d7ZSo1N2eXJdrEjkCJA/YNmM+0fPXa+t7Yoen4eu0SUiPjyJ2MruJ3Fg6nAejWzCVGay62mIpJ
rwmqIUeTONvghzmCKHbyBIxDU8lSg1x1Fmn1449FYMgkfZo98XEvXsa77hqtemgAylB5aoKhOlbN
Koh/lVckTvs+99drP9VDv5Jie1MEpWTg2ejSy103+DTB5zTV5FCYexNGBT55OAmgBxc1J8LYNiw9
kT/1PJ6duMxl/lo20NoC7tbz14XeFegg2jYUHh2sdVW7qanmGIHlVI1YOf106n1HWoltfCiCjudj
sSkKAcuFWnWnMIbvqRkDq+chFGhycOFIrcJZEbhhIzEIrRinbRqf9UH1E40aMLlcTTV7uoSVPi3z
PHwsXKfD8zBgChOXX1WS+v4BZKyvHJeXrJjfyVkPhnTH27B5neHznthA8f9jrQ50YEBywD2GeYt/
7kA8sLdyCXwxPRdFFf77JFAd2y9ppLlgflMRJyphT5mcWUdtPSFLzTy40/7+J0F25W2mxQdMZEk/
N8v5RfKsHKOQTrRoOnfwsisPPZSJRrOj0EeSUPFlqJfn295swgwGKpkRr0n02EAILrMWA2+UA0t2
UtJmdK0pthl+CdgPxWIP5RRRfjzoJe3V/aaf1Y9H7hkAqAYSk5j6DfqYCt0FwBA+udBOpso16LaU
3rlHD7mfk6rt6Sr54pZDYHb3bJcYwJsXNYbUjblFjwhPdEHqW7VdxNZF8LfiwyYSWlClvdcthoUt
EZgxTj1XCjWKeUDVNbjrGv0IiTX7/CQgO1f66qwmScJT1JaCrVC6DVQ/ASL7xV+Zclh2Z5tuZaHw
lghyIVKgQfGTpi6NfjZcRaBb+Iio8D2wmnd5xdxoEAwk2PofIi5iQNR2AsTdf9tcMG4c3N5KLDTR
eOWAXGbtveXGZLl+qL0CzOzCMjH9FxviDne1ycfNwv2iw7RZfBY8eTgtPgXZPmplDv7Ia0TvpmN1
l3/FIgvnIwmhYpyUN+AOK6+i6xpxXwqB86IcLMR830v3pxw6X/ZshbUHZNSMi6oZpNEKaKXAGorj
Y9W8IGbMFRS7aAP5s0vwnmYGVwgElkmlpKON32i5+4sjVgwjlA6u5gdsswuBnwaUgluNIIJ9YxcH
IbnR2t+rXquoPkRQP9ZMxRqkBQg2Eta/TUEj3o9RRLyFVCa3G3tgDVodlmRVp8xc3Nyw6mqa7hNl
IRtQ02W/cCeHzq99FNp1tu9W7R8LL90EMu/Lr3GvEzLD5cYf35J/ekXcRPEQdv6jPuMwgFLURysP
a+kpeA125n0TZobIGIn+tFgEEPLSsZpEyWjceeUrbDAOfvg0tBKbJRY/WHEm1oBQD6JBQsgKJ48F
7lctlmA+nTw53B3ulNRzUaPhfNgvUcLIt+kOP52YAdyaDBVzl4gitVDbxtQtaDEXFBwL7P30B9VN
ZUXIb7M4lJsZe7zRPzdpCZ7jOZjMlaE6A+/Xruyoq2hZqaHs1DMTwyQAs3JvyVpTsF9p1rHNcKs3
jdppxuPTsnqRfWqoEyL5C87Ok9JGnkYl9WbI5X+s89JfLx/ba764oy9ur8EIEXykSJR0fpkP6TLG
mhdoYBgR53/p0BKWa4JRwp5Ly5qM+AUlOWwFggBguTXzTNOCyW2ye1bdWN5wRXQ8QS9VlIQMAsIu
kM2OehpT0hy4FSsxcgUsikKbWwnZYaPR0cGeSE7r0+6U6I+RDS0cFRKpEZHfeFlmUW8hGoe7mL7F
AdaIbTQgNza9Y+M9vW6HGjBWO9MxQZMGa4vUSp36tqnzb3ijpU3BN4J3X5dDQv4+Wqiay5RXXlBa
xND+V1Mx3GzyN1TzJgrJnE5LE/YKcNeuk80P11hXgA/yFXAy7w5vNd9mIK3C6b0F/9RejEXug4ba
yTu8JwtWNjvupO1xBwWdz9JzF9HZuWeHiYUMawqx4CrSdpVOTcgMI7KaBbaycL5idvwLkF1/3xSm
COvXKEfZHJEJhCcygXBPXEkvx4DSpnwsjlEOdUdCCRG2/HyRQMMe8WgYk3eOLPuUAbIpftpE82aB
WVKB0PPggD7x9f1xPuO2eB5Lc0F4+4H/vir+YaCsckAeVzwHL7snhAQHmVvr1ibMoX4cLSaRTUTR
1tQ3cOBRG1BcdGc7z4JQv/t/ueKljIJ498xWxy9yim1u5PXGjjjXaQFIJ+S5wn65LT8EZR0GA6c4
UHNJ/x1uK4X5iSRvhZfvgvBZ3wb3L9LUY8SAic/B7X+e69LbIzweFmwllkQcWkKfZw2FIcQXdoRO
WgClCMf22sCN3/KSnFo7t6nYSMuW4d+mbNALQry6pBexXa3WIfo+uP3bRRYACsqtEZTvoKi2MfKu
O0hW4EZkvUre6iKMndatu5JVAsOATz5IYZKhkP7eBKrtXwiQP1G9x81zVgFubdG94cxgX4S+ktKS
iF7uF6lCnHvWtkA7zw62tk8Aqri2volcIGi+XqUXr6zQl+a180fK62JHecxslbaz+Rf3AgxPcIH5
U+YgPSfTuIJiHgLL3A+zzAQWoNQftyRKBOJCq/JUFWJyj9QYvmAk0nah0RXnMmH/hwZQ3VENrff4
4DUIf/+741qB9xsyWKO3nQi0ZNHtH85RFFtHA0N/VSWi/Ue53J1DnbZrXfqBgIrfybknuxOWeBXe
cU7tkPBsCXWuW1O7djE1sPcfLXvJpS0j4YAjD2Vl/AAjr1nnVXDREU9OSsbRK9Xk7qtV3J+0Jl8L
SIt2pSk4TSptvxGk7pAHQ3h8fLrCsm713/suTvU+s3r+lkXLIIFRXApP609fzWSkJEqfDBNN9zzY
a+8lc09vIeWAsg/GMW8KigRpPNT69Rklr6ImnpmmISZCk8mI5pSf3weDJ4sBg/tZMcZ9azNG1MKO
R2XDpekCcpGkoEsKZz5ERlkiExIwHvIHxboaeWYvvDTNs80NOP3u2xyFQvfkNNZ4LDLjf5eWTXgr
zlU9/sWWkmBQlxDibD8oOClXD8y9RVpTZyjWAIBShg7R7miymrM3Jxb5YWYvJE5/jdKWbemEmf2O
o+tvDGJkX7JEdhozAlRHq4WcjUl4NRY+TUCMO+XakBVzokbn3IetrsdPfXGDcnEVwlJaRiOsmJJg
UtQRu3bCx1umhRjhbUGnohniT9czBqx0mCRH2ocwATirgXEZkydKYXmZOwjCTKFW3EQ5HiZD2Czu
gAE8inwB6gM05F9n0+mtAfYAf0GwrnNE7vx7YPNV08ZcQwWwmKGGUojeCIDSJwBXIcgnfCLAqHhN
jCScw1BP1FIH266dG5kDVv5rHisOMfa6UgmIDlUoUK2QlI2+tHTvxP5yvYnkE/ucMfaG3t8VMWNl
dsQOTmr+e51M8KRYFmJ95QzlbrJMIhzDxDZ4IPQY6gttZ9LaOVyj9VzfQ88iVVRJOhZ3+mBMbLkf
jHGOg1B8Aa9wP79DJgwBM7DdqXVZ5+cKlpCJ8AR8v/S06dZTTp0ljzed4Cz0TZEpbTvbyt8pH9Lv
swIhT/mI0m6I9vBy2tUuqeIDiHXvIj483Qkg6R5kDHcCcE76n/074E9y7QLhZ/QXQ9WjH90cPWvq
L3ZZZoKhs4Bs9wHDMiK1eLA933HoYG7xNjxfRhY/jl/VZrUqqZ8mJw57T8LhQieXMVN3haKl3mCT
E7BYSvapc/k4m9AunOkZFW8YIeIM35LqEuswR/mFFPsli0il/98tMP+GbGMxHV2AjiTcBPfQtNET
QoIbfe2pywkWdL6uz6i0/cRdh10TC21+JAe+cY/BjUIY0pT8ijcHBOFKmSc8kbCPwspmcpETbd+O
WrYshWW4Uvcxlxn+lYBiIFz1ypfIspaKr1M0ZeO2WJccnW73L5UiXlmMzOMfuKJVgmfNMXKKuxr/
vjgwPyzipf/OtzDhSZ+0MisNPi5oor6O28IiJ2eLW0qmOEszdtkN4iEQSrm931TSBRmswtyU/E9M
kB0D51fRvuSt4m2qcWkHajFRwsdiW3W4XP0KwNW5CWfyq/ty5/z6P7oCN6O8mtpDmzybWk+2UUJO
S9CVjfKuRPW8WuTIbfoPMCAPaOyLTDQy3XfLMp/SVXX2A+bObVd4os2l0PBZUzKI/KjBUE5Oc4I8
k9QQ+2DP92d6kkf/DhHTNrzzKlSWy99NhpI7nJcPDkLssh+SsXkiBQsuWkJVmx/uPy6l4J6jkplt
hGeajuBcHo9rCtGuSn8AjQfUmdQoud4UfyikUpcNVmM6I4GiTn80lQTG6TxDe+mKg/37EBnc4Bas
jl+fwFln19sPxr9//8kNhIw3MANnkS3vG/SyzQrrlaBrLhyOzM9Tg/y8NQen8NpeWFkAQyx0jNV7
NPK0KTEgByrUV7kjaCxTv49oAFUpMx/okmR/VPF1M9kY2jFWCsTt9Ox2DL1ckHcDP2o1xeIp5ozH
I9Etol5V+mE1wWlj4iQmUmz55cTRlk5epVOhgrCMfFpHodpjMJFuWIthrTv908A6aTx4vI9YQRHc
gPu9mKOs/SRx2FSxHWiADm+XFsVWpqfWE1Y/IE7azf4Zped05OXPnifJ0T9IXlcWXhTj3AfHRWwH
SqxrwJ65FVuO+IpAj1ctNdQYy+lbwfEigy8Vdqs+H37Qoz/RMY/yEYN8bPF9DjmJUGGBLCrFlfYJ
k3DXDPhf4io+Idaxiaiua50ImX/4F/RyvMs87fstZIINyFsH6mYa717sAYrgHTU+kdKWU7JxGXv7
Q4T4KH0fMDKV/Ge9Y1Li5J93bCPLwnOXplHCcyrWHKnsEE+BIn2d/DcnzMGP7dOHp5mQZwEcDgj0
qbcx/54hNCZEiOAXjBVKUt/xBFbAlcykQ4rDQUQkeWKBIFhFCftSIq1PsN0APzhEIV8PWSDzD3+C
C5xfozHANSourY0MSloFod9nDfP0SAOP6JwlyOYZSF8Ftr6H2MmSkARIF0b6EPQdDH46frcvr78T
RSY32GPuJ2UnahZetTpTETM1OyEPJVSCfuUW4FZ9Ptojyrg4U5ynMkYNc7Ebf/0noD1SxZkJVNg/
Ydhz4Vo71r95rdbYSj0YfdXCE+RwRFxK7pA6Qd06TpORygykzkEhL2C32jEaHwXCOopMBjIu6lma
G2Z92VEtwxcUiGM/eEtv7HdiMdb3O6qgyqT+/2wv0T3pnZl5fpXOdtpsXa33B5dA1g0ShozBl6Cj
MXfggsMIV2r7gmYH1yb56Pb+vtG2hY0R+icV+dK2IgpglkwqKa11AF+Th/Rr4VzrJZ8T4CQ8gy1d
cx9A7Fs0Eq/ppUOPCFt9i5m6g5EzPoamR0gC8HlaDF6Z5FBy1BMWNxFy5X3G1DYseaP3VV8Emjpd
lgA1Jh4KrzDLzF9BPnBgSQw/S9ffAr+lIZAZNktFhgXnuvY1UrVCksFNZiIEaOy7/IJQuti87m1h
b15aEWMeY6mLTJnP4H88ARCiJigCKgnDN8br29Rp3Nw6Cfke1IJh8io/sX3wPVsZ/dyQCS1CXBcC
rJpsK1cn3CrwFG9R8PfDQxYsKPU3zgUH9ms72O0JtMeOduNOMxxWLpcYrxbPpvugCII1LSc73tv3
svagdcx4+dLn/FQS0EcfI5X3wFrn3qI8+e4LSn9QtqxBPiWB2aZ+B/i23eM9M9aqPw4Sq7hPvH5z
qa7DXFe/5pNwvQZ4BOoZr8MBQ3Ii7AFM4r6R5rBm/TYSf7SfAVZfa5jBwWMAgh82lmFr7BG6byf0
8UbHZYOsf0SKEqkCvxUDPkVWr69zHzGBYuydXBL9S+/3WwCP9B+6hiQO7jJgz88g1tyQMAtVwWNd
Td0ImBLvNBUHTbriYE2niklivS6uykB8TA+vVYTXupZDseXYbnZNlGEnN8hiWmVE/nmPdtiC2IdY
PipmFbxPUVX4UJfCeCeMYIqLiWtcsS2sssQ5QHRS/Hz0CHS8hlqdbtVCV1OUquw6yaccEk3vkIBv
hNerAj8vNeBOYvDn0M9hu4wBVkpyH9SlM2ugHxeB/oHNjjvWI7EZ14e5kBUcaZP//GNJD5tkr9Sd
2EPJZqerONUYARWfmPwogfoRPLCza8ycc5fhr0oO5BP3mqlzQUi6X8q745a7pUrXj5vPp/pmBALt
7dpYXidOjQuGtdHcSk/jX+utIuPNMu6ouWYOxaV1yc7TBBxLeo0MhPQdt8GTCopjH5tXfvF8VFzc
ik6ZNQA5FlX1yM6Wk2ClX3IrRGMdDqScXGQx9f+hYP4iAGB+pc2/aXvQ8jhA0sY1Zknx1S65WlFA
SRSuuHjbNRFeh2ezDj37HX1IwM4RzXJ6KfuG0E+np0h7XdNMTmxoL/prvfxyfNsLcRRr5Bbio1L3
WrLe3B+9UH3PDwOo3KIpFVD94Pz9GiWVdcBqo5cSwl4EW0S5fv5xHchNWQ5KHrgOB7kq3e21m8IM
tZ1/UTaz0epB2kMRQ4QlWDi9XrkziEE3GdeCAr0EIeK1OHQ/g6zl0hHJokLXxB60BEyUBWPTldlQ
Pd652dugC2AIcRk78pIlTBGZK7EFm/Y1Ppn4BumqpGOxhPH/yUk7FyF1U8iQLwYNFi8MLE4sbu5x
1YEnUIYwbSo/Tc/VWC3BFT5d1rwEWalwIPmmeyRFPz2+D+BI9XgTCUCVQjp2S6TFvV9m75juju9r
4k5zO93JAzfxYVy4G1HEFucvFeEVBPj4gy/sqWqunfRfRZkgXY+n8cTL8M9ypeLsEz0w3ivbpFM5
TBeBO/jJ/87H6cr0U2r3glob3M+na/kZ3bIEX240goHE57FqjCE8s5KGQS72GADbRw7lDqjxyNRE
daDXu2ELedm2x2IyOC8rtLKAwfQUCA57WsKsho3whSf0VgCaENGVGBscqNSSOFZyjlDtjBlYadMF
IM1JRye1ALsNOMwdXMcCOGQib5NXkyz4B85ZcKYZJUo6/hSqrU1y0e8oXPj1sIRWEZ5XSh7eV2fd
0CHztyg7N50bwE4bAp3pvWrZGzFgdWOxIOtp1+3kSWnKDO8eFR/y1Fq5EBM9kEpVDgOfnEITDZ0n
1ZrrX465Xb7vAY1jy36p/+/d2Ctb5ZtaxWpIG90bIfHIZFiUS4A9K1U7K3sbzJSfj/XUk45Wo6uN
8JrEsdNe68gmND2lTUspOoEPw4PKjGxiTB+fJB2hePac0eoZZf9o6TOqrv9ScCfI1I9k+Xa2uSWd
EaVg0crvDBKXKR6U4zD49FDWKl1RMTz3xAiSZdwBeCDZO5rv6MwRjPDGIXQmPxT6eIyg/36qAPtM
pF2ttLW8xpxzp+cW3d3dl+oTTNZpfm9kGKrje0SKYGPJofwif2/me0b6AeUCgdT1/j5uMpoL2vaI
TF2CYLFfkK9CuWkMM1fZSFUtWRlbsETNo3zdVH38b573dtn/fCmr2psH/X/ITALa+rj08hg1PqEh
ool9o0F3QB/ep+BwbpHT0XphPp+Gy0GVXTjy+E/wjUs3rFdYNFVUn36AI/TaHuREYHD83vofIeIv
kddtOfx0OW5BDPqxVV4xn/73ux0oA5VocAjDszOaiWb4LQRGoTcXo2zPkFIYXgKIL5XFOGvTVJyA
ssbRQl4zdCa/JNG20QPyzcoeXttmMXGYIAnrbLvqalBzyqu2ESQCFOdIF14I6RTMe9nJcspkzc/V
YnJm5B7SLc8QM6PPLCNwFFDcWVOkoh8neYiv3ZlxzOpy95OWTaU18E2FnjsrA135bRdh4FsVBpNa
WCyg+9X71HqXAv1BFdqsqkXQDpwwKJqc2JP1C5cA8Cqs0tNlqObpgQG2WvbDhExq6/S+RRnE12xQ
p1z4c2sIW1HIqqxpYWi4XXmfd5TXmnXKCW7tvcBW5yeXZsHd/K5MdDIVUo50YkRf5AGrNMYsasJh
b2rhd4AqmXvZmqz0RqWNcvVFHegyy3SdKgvjM7lGcPlwVFK3Ity4Rjbt2sKW9htiodgV8rbCq0mA
2PoUoxeDKCgvIkIb5RjvtrPtbGDKu9ckY1+d4c+47PUdQul1dLQJReqo7WajzZScklmjvmirkk5G
G9d4kFiWrLdwBEcS8vSJRITtEOrk2Z8MUGMekAcUuD45314K2t3vi9mMXU5LaGl5CWAfRHiDBu8U
EJe/1R3GcIhFOU5IdMtlMfkOmqum1QRyt+EgjBDAav/rueI1IUBgDVDXpZn4DOqCiXhL+DWaJhPP
U1RJpFrAf31jM/37cxLxuopyCYzjXRk5AMeuJ16AOVn3igVcNXCorV2Z51bfvKGeMtkcFaoNroDs
PqoJCWSac/dzefmFoU3h9Vs41ho4BNoZz/g9FQVW6MIwOaIjrb42rAZGcpSOVrw8Upo03JM5nE13
TGVaH/AeLPblBml5H3NH2ahGAkSiRza9nSFb2gM7fs9QGBbknxohjbf0uEcsUJMcuJ2zoJPAJlw+
K38isL/aYxbFrEEE9uZV5pR4N26xGQT2v9cQ8SYNntLTKgm9cfqWltytJbW6EGxuP/eqsu5bCube
oARAPZ+EIspuFBT+/Qi/fyGNcbA0JumXiqoWXy+NL6yKEUVf8HsCNp+cFBToAgu+0eXZ3YdbsXRy
WYsscK1QLyxsF4Mu3Gh+kpwcq5T4w7iqHbvX5m/f/PFuBKlFwOj4RQ/a08fnlHT5V69MK9YAM2Fk
IsjtrEHN7zW0CyUm4e/ml9q2LmIe2QnNyVcAAKUQSPenQXNcyLi7LthHrIOsdF+oelC7x8mhTaeT
6vka9Ks3KW5HMYSX6g0MJbIim0pYZrOe6KGmbSy4+3S6wS4dIcDSayF1ZZnwuVXbDienlx9+P9HF
+i3C51f0YygDpV4a5aOUmH8NtYkljNIN+6jVvvFnSPFEqN4QjmiZS1HVEQY0P2j9BnPTMIPehjoH
oG+bYiKWQBR+wDnGuv0ikv+enmKO7sdba1PcJYUFpFM7VMhOMoHaQ5B5dU6U0EkGS4EvLcZiuFqK
ezoWEvUjL7A+e0xaRQ1omgQuCPwEry4I8VuREqY3RRKVMpLZRKGdSJwCJKER6r6SDEoBi1lvgY/X
JlUX87fC2SdpYBcXm2f1MHNP6CpnMQu5H75O3K6DrVX4N+jyatRcm8QMToElpvfapALu/6idrFvq
YJE7NMhYzEylZLtdJPnAaH0Vqar9qbeIcbYWC1m20FxkbtjfLHjUzbG0DyOK9JaDR9af/879jntF
+TBisM0zYOp5A+a09sxLj+U3bgzCwuzaWN4sE1YHFFrtaRz1vIjcPpkHpQMwJgigs76TbATmVTfv
ebVV3YzyiE3uNfGN4RIZc6vRKfXsbLS97xsj21ao0VrMQ3sIimglyLa2LQscYavBcX3eEAzz3Maq
RDUXfVHfthTCphi0Et+ccmhfYyobMZDZTXONH1OF7qVF23Iq8Fl0xHJCbHdJMtoSzZqk0sb9e2j1
RxljNFmN7sRRSC/8wrI0jgb5T3qQJCACCmcdz5oxH9jQjX0SI1rlkQS485S13PumpLSLYYKelcTU
6wr0GzzEHb7bNYsZBzab4DAwDFMIhK3vvNVLB+301QTt8ODZb3qHwYFu/RuVrbTPInwvx8890p2C
qiFDgJLSaOKHO2DOmecZPvoEF2SW72uhh8RNNzdHGy5R49jnpey+Tx5eihNZRbut5249eRLp2C7H
ygP0cbaZdBv6hubegoZoVZ9C9dfUhQ9O2IrR1zXeC0ISqYkvW8m7/Ke5av2c4CMEWVAdFcx+ad6v
4SoIYl77UkEdhLNjc2yr98Sln0PYjh6NYTFyTFd7+7u/RRNiYhjfKrcMse2xXjPUrcwLLIMkJExE
83BsaNPsJFkayGrXF2oYyGb1voXm83DDOzUyf4ZBIgjox/TPz3rduYBjDjhIGVqhM8v1YNkZOQYC
H8MTgPkxgESVSjma66NW7bhkugnqeYGicssMvWsnE3dhcz2w3ExMJOYdQshdxoMDQs7Y0GDhy4HG
HKNL181kBW9nZP+e9+ztwB+15yQqVViHM1FxkB0pv7iJDR7EaYP8jMGXVmlsioS8HnTsxUNW9yDz
PkUT+0YhbwBfB4sWZe7lbnLvLaGlLxHnu3yAWn30pWST29kuS16svZCrNF4AJON5AHPzOH/wp/cT
NO6Yd/eMqPe2bTJaIzhvK0/TdCYdBX+um9Kyi3O0+4HGovvCcNhNo7kANq/thgPgGJoqmipoIg1V
/x/xlgxomK2hWylxr5BZw+gsoMA7yEahODujgroYZLKD+iZpFMpLHZwZGB2dK92485uRW2ZLCcWn
/1Jn+anXOo+krfL2Wt3mILmX1wYZuovcJU64bsmSxasQ2d+OK4QlmZBhfv9OtsYWS9/oDfM1fXKC
onEvD2poPSJvQrEEFkUhhaW/vOcilj4t73WxcySbRZRDQFNa42/E5dQolffeKABdKkledb+Fga+0
fWKPDYBe+YmxGUmXrBE3uMrSAvVgHpHMICgHNcxnzgxhlH10S6m5aquOjUGYm9a2I9zY9ncbA1es
/m6+ILIizGFtVB8j/aJWTttOsbJTUmBKlBPw/eyyfr3omTeqgsX2ZfWbNOIM2AquvneixxwJ66+0
eRbX1myK3abGImLcOMTRGUeQ8eNTAS22ovreOq7yNfhTtMD2pOVHglBhRu31mTJlqsJOxxtuwbLV
xOHSYW5YMDmxfBuKy8vk3AXP7KIZ9cjDm2FpuR5UlK60sJZCnX02sK4i3kMPTsrnpqS7lptDHKSi
+XnFjyOZ2Lm4E+g1r1LwweCC3TtXzPu5evCHmHZQWjKWdsh+BkbEqYr1XwMhG6vXiRfn842eIfSR
RodCEvLTIWY+4TWyITKQoC+zID/i5h6RiFtYt1CafNZ8rX2B6oniKCNyOBmjEA8jUAqcsqOdaXWU
TphwBmT7/cW2Vrg5uVA58eH1hbPDWBFmly18LIYdC0AqSq2NT3ucjLzoYZCs0+X1Af0pD/gBk8l/
LQko6Yff1bzm+3gXrBn+Zm+WGo+GcPrAu3p8wbG6WwbLEntME7VA31LrrUXzIlVKGyKFUyRGdBHl
ePmpcLQ9xMK05hJAQ4DOojD2XndWTF7fJIaIptJipmPILifuQ1nFlcX+YWJzIeVwfyiDBuNDEkWx
KBUa2ISlDPLkL2/UlZSHLomzNhC686O7LOZ87SZB9O3ylRm7qolT3rBYTPfgfBx5JepGsVi+mQEY
iaZWEHzNzYi6P9O3WxpRGdk+Pr7mGpxSM3GShaP90525Xbj86TvumWY+PqUJqvqpnhESmwb2g1rQ
MHTvFRjR9r3em+j5ugPKjvfpf4xGUL2UjYol2usC04Wmsm4nRvX+qc/g1Au37vx/JCgQ4WTUyhZC
5UAkUvjcKAtE32N9ziSov5KIOSqR6klONsKJUOihOslHvFn8LwKC6XGLfKzEFch1QywYaeRRk8Vk
42kktLm7fIl0jD0r2tIYRxgMlCuCdx6lClM+V0fpSvCituc67MdwaPoPVpyF2bKJOGVF7coEADJA
lv7e1SyOHKkuZShdV/ADs9B2Dkz/BQrteDSZCoua8157mep/v4da3ZzK/ppNarxf9jYKndpyg+JO
jH4b/Sn7Sbl5bmDxQij2hyXb3OxOA9xwhmIX97vWEcxKSoZbu1te6o+6KLNYbyrEX9Ns8gqf9sZc
GGTHcxKWg57kCiZRFqUDnDq577KnAFAnlExg+H4SeSWMzojPUjVF3sg1ZzgCoW3LoS9fIm8Ja5cT
vyARb/kLPGuXuagE7Jx9M3KkOJrS1p7a+4c+8A7GGEEn2XLRLNpzmF+HP0rFk09HBtN1d8jxtCnE
AK/929Z+HhUpY4e4Pl18KkPk9u2831i20piXqQt52wFefmAMVYcCqTl4s3DGrNRe44fpdtk5rTvo
2T234qMRQ2OLZUG1itES/MsqgAOCPifdFbYZ0pHfPXr9lMYEr51/ydxahM69gaALB+eLEHrQF6xv
4pzdUfXRPz3n8ok8C8eSEME++z4YNaE5IG5ihAPWy3dREZ4IHkxXEv78Ygpd4lJA6tS8wBJiwN3R
umknXckaOhsLRuWftJaE8SWikh29kRW9nvxMRQKMY5s86q/c9pzR9OO4QQuwVCwk1N30sUnpCuZC
ww6TlSZuq6KBRfNNl/+lDJIl1d1ua1VgLOdqJL/HjuFqwMsXYwONEzOIknxG71uv8hCwDQ49YoW8
+MYR0GsWWSb+Q47Vh4eBWY38V9t2PJ1mf5hQ9HH9t/wnCgfDpROmcALVL+s9WBnKvcAJNBkPwm26
nUB+fBGOLFW4EgQf07xfAS5uldat8bleaiXp74/wzHkQSKkM3Sw/zumHd/eoI4WsyonZHmCyJ9Qn
Em3yOulnUCrS9lUsLQHwa9Ox6TJxIcoOzhD45qE6qnhkpfyT+5YIT2m1dvIfgZq5W4mli1iaB6v8
2e0RfsqTtTxloAwzlgzQ0pVVnLWu/ntlW1Fe466A4cgfDWYAb0fYOMJqsAchS+JkKC1nNcB1uFnM
gNluQ33h6ZJRibadm1qk0NPpMrqThylHARR0PXidWDQAEj5iY53RD6ecMI/2zKOxhkINI1kzkqpF
HMwyxuBqPswMhvXjFKg0vSVubyvTyMVBkFF6YgYHoF/qDTe5+rIgF9i/gYF+aSOdekaLko+4bJZj
dQFRgcTTqn6fC+2qUC1tGW+bNabuJnXSQW5OOYf9xK/zXHkiu9FsvqwhCD7RumDwXY61gR36tVcj
ZbROnNe+RvR256jmc4nXlXJmwf2CLjEvQtfBJp/WGli6bUwSMRJu1iBUaK17vIzWrJLRR6QtYkPZ
I5aZxAbRyxkq29CylvWCptO059oDhyzVqzLSsNWVYr9235sCbdnKEoPbiJFuP1CEyQN/rZRioW5L
oyoBdf2pZhKeMSNTYjm27XSd/nMQ59X6wrqCUKp11pIMAGswpQAw5o/BVL4EJvppwHiZ5s3Rmepk
ITzeG6Zk9SB159S04c3BtxssWcfRNaPfIslmsGAduwEZQjQ0age8n1KTpaTSHVDEmARXckrAMeNV
Ry1u+v2Gt6diulYWBV8Vibzxih/WK/QdS5F4LE/SfZ66nqo9NNrGMoYLaHu2RmOI6P5j46RCfHNG
oyCo/sf0swpU25So/kgU/cwZvphgG7Swoq787qB+U1hKquitsyMgRhX1aUGYO+dWH1MnjWKT3pya
iNYTeNh0g4UAlUQfbVZbswOLbwW273RcD64C1zKTkeauH1v3smWJU0zc9cQ/HNAo2IqbIm5vxkY3
OkIb/DPKR6D7DfMkRG84b1hchI/dmmaNmkYMoDYwY2ORUU7XO64h/SZLEG/k0uncayxrBP284fW6
yETnIRETBHMCCLBC/wmqaJpxmNTpAIY3SUXGXMH7kxGq+siLqTi31V1Vx23OEMShxIOKl4rg5dUO
i2VXekOp2GdX24iWJ/csMC417XCrC4FyGRzn0GD4n5whaUhImjhsXZd3xA8H0BkmUhpc7BMndpMv
LIYYrogdxQYmhbUN604YFgdfX1/lbiHvgQ84Fw1nRWTWygqw52oRdDZ+V/05xtrZewhIRSqqbMuF
LnnIQqhdlV3GZJJdzCHEegCQvb2iwhQaYgA3KJAoHD9FJw57e594II2t/s3+J8J4RPFeF90pT581
Emq1tQG8eeuIL5zaSnfk49/XndegYtLJfxSV8M2ZaDMfrHYXt1HrE7NKe8H72wPK0QbAPCb7CFZn
cPkmGCzg41G1znayOZ6xxPulKRegvGZlluL0t+ojXXLi/ZcxGT4UqoBr9UiioVj6uNzP47ZDVMrZ
gYfN7WEJrM+eTEWNFtzQx0GZD6WsTYIrUsBo34kITlhR7Nfh/PaG/JqZCIgOHAqIJYdl8JffcHEY
YO9vfAAugMuj2JsWuB19dpViSm/x6ADQ+193IGVOhDoEdEHugxVMPDuhDKlDgwDomXLtC2slJKZ1
qwXN5rOtzW4ZcSs8+YCFIdtf7nGlwP5aHKgYwtikhnRJBkwrO8o2X5xPCmqpYyyWCQpoCdOzBo15
qnhD764PbQgadZWNpwVFcz/YOvipnJEmyyhAYUV5k4Vftf8Kndyz7e/Z80r6llZf3Jf9OtVTNqTG
aN5zefNxg3AYX5HPQQVj+DNlcEnkTpUzMPXhwnUA8KJyt8Y72OINRPZPTy7S/AM1rL1YQLMjZbeq
L2UsJmG4ASs6Gih4yvmYrZEyxqWNTHVCBqxouyrCdWQIgFG8G4suED8eizyVKc+ljHwrNrN9WvSy
U3DfRH+E4dzOKNVPDqbFafZ6xJQSFnr4GOGoJHIb3uAe8FDh0x4fvZW40EEO5EoDKv323hFGY0p2
3/dBJpU6Tft7Zk2FBMarX4ueEB1liMG2EQxceNPEY5FHMXuY8rlwk0Cl7/EAWViV3utI82zi5g1L
CpH73Mq5tsiSjyE9onhBMuhiEFyuKys7KTOKLaZ5UTDe9vJOnLwt/tswvgegc7EoIhVeyeCwt+Zx
s47Fme3ABzZJdrFrs4ZcAiLQa086cnmM9qo8rTtkF+0bCly8qO2dfdbPi9qnznjTEXeZsvyJNI94
KkEI5UE0fhis984UE3FqdNN6JofK+JJsTN56tH7X7qNBV6UXbSUoVN6b3XHHAdsuuv1AfKGt8DNN
3IdZMeC/Hjiol41vSCWXqZVUtNrDtRRuMtzd2IIS3OB4P9uvlNVWvlpARv2TEP5b2MSyGG/ux8et
C7LgDHefj4ub9EEWW/ijUzjksq8J4rNhNjZ26ES1O3R+fy5Dt47A97xd4OSlzkacLt7Em5kWXGB/
4zgic+YCH5ngFZSBAjjG6aiX0ECmV4B4FI53KgQVq7lsDzZcjlhzHHhOwymXrBK3smqYvlkrrI4q
qe/utyBGdfGRXJ+bxIAMKNUIFF3mE/NnGO+n6kiUy4hYx38xqubNucAqpBMvINnfRcHfhwq+m3fv
pnFcLZ7un4995dLWirYOlkgV28In7H1gDsmnhvKT94ZNSbu+wb4a8N7A5FnbOELVp/PrBFrtnff/
V5Ri6XQrQEYEXu9ZgoTLY4ecoe+rMA77GmtOmvdUNhIOxItAxIKEDYV0ytMMrkqiuCtcI/HhIuxc
rb/LKSj3UuhPcqdk6bae2jo8L1B/zFTmT91Ok8wykFxFtlgwE8xpbCD17CUU8sDGnFSkmOMV60HW
+ZLHrEroTE3jevJWJKNyb9VypAZYjLL/zn0PjC4gjmmXEe9I6AaLOiDHADpNfebyRKgoAVBPT8sk
jwJNmbn7rLQW43rqOZupsJM2J22x4fKhstp5kNQuT5FANWxDd9o2F6KrZ2XfZcMD/GSRXVnkzRJz
loO+LBIQ0WzlLqvQT/GSBYn/RoZ6uXQeEW8Z5xUHbDwIrI/a/9VWNi588QRoLnpyiPZRb+6ASvjK
0gSLDFB8ockmZ26V6f5fPFwwgsL9s+1j6EGWwLfL9RzvcpDeYXWE4ZtHBg8BnsHSlwlcJf25wklv
aEPWRHxR6ZwfVOqqSfHnKDFYKLqfA94ZPTs/fLfnLZC5BfxRTcF4Kphx4R6P783M6yX6OUX2amiM
mSIN46PuYjcQOI6AvyslKptbR6lUXtS+PRvmMV/9q3gkGYOW1ibSoVs0MsLFZuKQB6E4r2D/pcSp
jXngLX5DVWzWDB59v+R7wvdTKCE62sTJMCElnsL119sOp+yxU13TkKWAQzxZNGEUQTHp3DQ8cXLB
i9n4vlqYR6aP9JOKU12N/TpP2FFSsQmyiXy8bTH5y9b3EJgD2tBcIPwpu0GP5pf9xHPWOz39nR4Z
SGO/EOmakQ1YQcie+vfqV/O5zBaM9r3Qm5vbBOnznjtt0bSN5OltdinJHNFGrZfyWri3ETmNnI9R
joCBwkSQ/fX89so7iGOS07ajPoR4IDVoytKTlS1ouCRjS8Y2psYDZ9iKY7mOOR5e6WNAoduC4W9M
Z0YCELQyw9aqVN41KV/D72NGogMIrpx+OKLZdFFDL3jYuNWorSBYmZdHVi33AS3tmNC/WsQRHoeJ
xWXE1CEWFvgqUVpNcYOreft/uFno1ip/gV5ablO/zvYjA1wwv7z8R4rrx89HTr1r8K+SS8409vO6
CGKSqYPUWhEBZtq8FkNdXsH9GVG43lvy22NBpkUhcXJy07QGUmTj7vf2TyBqfRjojtyF7DPRXUav
hK5SUgxf1rn957NToo7Rx2MOk+U8ncceVatcwF1rDcpuiGoPjUaD1EkRLbagQKCEcqZMvT0Q9iMa
q8hJwuHhpFnh1R3G0kVznco+nqQUe6qrCeQ20mi41dp7Yc4UuSJd9WG86PeAucvyw9Qjey+nOrxk
C1zTGOK+/nReAPX2zGTX7YggkPr6aR5rdhevfBBZ2PCBPghZoVT7pvk52YlkJyBYHuG+KV9spi+R
RjDj6rm+rAT24xy1W5lFqNSyx4oI/QSS/sSS9kP2Tb+7yvYkTBiimfsWf5PLKi9/OWppEsu55KHc
PAVF6UX1bQuw+AN21Bba1mJOapZrm9WRUOIyhNF2+NwWEiuv1B7pVo3wBKY33dNozmE53IOEvjli
R0i8lI/LOTGNyjcic7LCMl8HBl5jEAk3SFp+rs/Hk84p3RECK2qZk8686Xz+uCWhhCfrPnBSyy17
eOFtgHpU3Kx+xbxjXhId2pv79HVwQFLUtdVc2RzpYy2AAfKnurhpGVRigAkU+Tu49PG/0LFNoQ4/
bYF9M88nyudVODMlMfhbbt995tIVMKoVJse5fPdmFdCCPc0ilREnkzHcjjYcO0DtX8hLf+GFlMVB
H8Pev4pyBLSS68WpVc2FJA+86NxCaqqWwp2ApJ2pCak4lnacijoVa4HbkFecLBrJrt6KueqMdPzN
LmFAcioOSwX7tEMdfSonaoT+pjmfo+N5DT0/7UsrMlx6HZlISqyQceeX5oBs39Dal26aNGaUrkoY
EpcTwENZ4u96YX5pAdjlIzfxsDVCCpsGBatxm8GnGu0AfWhp4zKbtW6NPXUvxhwvDuLFNX8472yv
zxvRWozWFZKl0yAgR01PiUOPzcBTJXF2ZUrhkN04kDSk2b+6ZfXurHnorrxRRFPMOumc+Gmq0bZz
7OfyJAyPmzBcU8ENTyh4sd+reAHors6wexD7RWcfli4cuSAHl2AWVwYegovzziRszEsRs7vceUaK
/V0baFH+JqFecW3505HJT/DG20SGV5lWFpVXEyeTtDw38u2TDxTi6z8yFApRZ5f53JjvRxiNrZou
8sg3r3VMZ9LJljmbfuVAf/fSAjT4PFmHAyg9ZZWft/UlDQHcCowcw2RCqJQjRYCxG0sII1hhpFUM
+HUIWSUgBo0gytbIOelNCDbRsWHPmVZtYqNwHe6OjBqk+1Nf+Mzsn6sg607EJpRSCzPJOvgq3x3H
nZcunUQNWHYSsNVr0HwDr7qA9A0lxZ6ynRnoE5Ag1t+99+OTnyI7mjsxMfUtaTjo3VydoDuFuwbV
xuvR9mbYTsAaxqXEbsy3VUOEG+qfSVdn+wchlyGTy89nE+GmsoqUZRR94r3QgK05NbvV62IoiJHf
LzSQbVBfTCy2yoDRfKA8hGauaPy7oVvTHuA2BVpKRqE/MfUIP12qLFdrSpCMoM8oLz2Al6WTonKg
eb8chmK2ShhxrBKs4lnytkKA4NQf6YCVH+Llxsi2vPqkJ7AT0s8Zv1iOtfa59oqXNB9JR06eOY5L
P8r3eRf3f06kZftDea+Cw+KKABwTUFAvlmewbMOIAMDPqPL59UTB0RvEMW6AKarqILKs8ZQDuAQ4
zT97dkQ+Sjz9w4pYp9p5WjO39nMrV7O8gQH3AWYAaMDADmRViAua/38X44VnD4X2n0EeoL1WfZu5
/NMrFrzmCB9+t7RuAVFhmO2s6HVqwVAlouuvxOkgrY2HdzxpWx6hAaMLD6ut0qfgCmCrnq/dJD5e
n/L4YQfjo0o6mS2vNWJDiD0wwV61AHgc4L3KfcrL8sHiiZC1f0R0g6bUfSFZbC7dlOZW+JJoLTjl
k+8LjEJhI3XHwhFMW3PcBZVS0yv5nZi14CzJgH6tvYxJOjXKQ9dXzGuSblcVsAPRd+T7r1d9Znht
pg0S1ozbVUBOkFO3oDGBzDioG4U7rlrZ6uH6er6Z1Mr+afW8l+zLG4iEmMUg08V9Tm2Lw5FbRczl
2SmYMcroN9wI51wl16qIQnWQRWeJbBJznzExGeGSe4sdfyAT5V2L/hZ7Wx0c8SwhJWpJlYBd/EBk
IgD6cOKwi2N1bNKN6veAcDk/1wfDy/CozvNZgqcdNWehEbc2ORJglA49cHG2Yxvs9w/YtPkcf1KV
KO7GaGqt1vvl+vO6bxFqXMkMMlSR3vy8mPnj6W9eh4xctvg8vuG+Xq82etuuEZaPjlzPqd0B+WOs
ipX69u0Uvt42o7k0DrDLsUNCbB9QPyntCUc00wQ3NEbNSgtwp8grlV21JZH5x5pjLBTbKAc/xW8O
+TuiODAC6sPZyxLmkyyBZ0lc56giXWJfpCFJRmL19/LrGFmnlHZsiDcOG6c9ifyCXj2ODBhkz5/t
5cPH43BYdNGS63aNbQiTJMj3fdZ3OvECoI0z5A/HeNHyTzuT9tWM3J4vg4ihpar2+V/MpubzXG88
OdhBOn7oonrjCripp1q2iOIjndPUDSbWkkiSpQjdtDvObu/jVO3OST8Wsd/CPEQd4v/r+qW6/MkO
yPF+kLb2gTeSF8x+9J1lBBOiCYacmo2NkAcrFHtVbpoVHqEpo0z7m+m5aUL/MhF69dqmAUc4KNaz
xP1tgarkhCgdGoCM2Jcssy6p0Z6iM7aSiOCrKeqKHc/Bv6eRPMCqOtS0e784hgKUpF/IHn1nS8vt
Bxuv8euBTb0cl1gFa8Z/SifKa1iwb3DSMbrXCkjoA/rRWfh2AyW5yfXjQUmoHJpxJh9e2XCel1WT
XnZ8cgBLtMCzCqCsJZzbSKFTLQiJewqS5/mQhGY5345CVHUw40vUEBGCnMAYb6HFCAosMl6XYDD+
kSu0pKr6UA8mT8DLwTXC5w7uxQSmKCah3lxjhfvkgWuIFvDlaPMA9rwf4AQsgfeVYLniZf47tftG
rqJ/eQIDhKEum/XFiXsGXWhbCwf4RBrr4vOQUG7WCqb9xhazQ3Zqe0LZGduu0VeyspAWd8pcqG0P
Uf0BGjPrNRBpIIT1VjxiRSlkz20ab2Oczba3i2EWvBQTeaLDSw/eXg83aZ0EubfllwMxc90YKjrp
HKZXnwLA2cKkg5c+m7bqfqqqLj00c7L+VMGoltk1CMcG40DV0x3thqjvIoObucmSxdBQJppfP38b
pqQSs6JvpdXtY3KDpfTQ+Wt2Ev72OSXNyV9CitBYdj8+lwz4yoev11OfhvtTFxzsOXaVGLs7IVil
aUax0qEeUyAiYaO/QN6ugPhWs3kR/qfq/iXB93Ia5mpDlkueC3Fv75m+N80HdzNdqMgrTfIwRHEU
95G1Mj8utaJGi22FkgHqos/SzqeezPMmlFKVHoITr9O0ogPeu8SUVnC7NmEJzyU7mb1RQkuUgjGy
hwX4Zi6iYkil2EfK0svKkQj12IAeJQ0A5IxqCPZN8bawZL5jY3qsbuR6KPKdvE+LPfiEk3su3bcI
gliTrQFhGSzOHgf/j3HMsnvPSxGSDHCK5cAKYk+tUO2H9ekne7B/j+lV+vdGVWA+deEPmwuCJ5jb
QiYaroMscNovZqNGKfihlR/6Esk+qCnxn929PAiHvBvB1/X1CwSX6zNOdeQR8qMSkf0gMBeYtOzC
OovilIySwNXTCMnEaGLodt0HdeS0qdWL5gDnyCRlCS4kIUkvgqcBA1BchRVg2ySekippFBnt53rH
JWyOSD8DRepR1uU40Ki7bcwPBVB7jGn3HO8JpZFazUzxOWJOKaLsD7Gl9Lgj49HecgEfC7WP6LOy
zGgLwjgrI7cBdHuWZ5dVIt0MT2ebjS4S3JBoyXE96OJFpPKilvc8orIwUwMc5nxEFHzpsMYA86Rr
DIl/Vwzosqk4q4+6RFV/bLa8wAKhtye7GyeS9+6EAjjR3NAgRPC3v4lI9W8uj6qgkHC9bUuvkUXE
C4PYyntgej9Sg1YXQO8o6am9vTYpWlY+YHAdpWzk0E+dYtg/tA3bdFCEz8w2XOVf/DEZ0ND3H387
Rik8peBujEyi+88bKWaPjS1bQC9Pb6tXqP8dO4Z/xl+UlasZT5/SbUQoiH5f3uIxH1CSlp0HzRI8
pfpzTxgmMcxie+CK9ORkQ8vOGsSK8jV/KyHW9JOUhp+8nl7Coy/7yUH4leCxoTdOzXjvjIoyPu60
ftX2o60kWz0ZjRLA3mizKPfTuE3qD9kp/cJonYeuUZrMdUZfo44dHK7nmtaSF/0q276Q3p7dmpk8
sm+GYCex1YUipvM8ggqrT71McHcsYOBDCfgH1btCCrxz4LoB+/JT5o1fuXAS4KqJBgiD6SVZCegF
zt8brLtm9Ib2AdvZzQuHg5U/+tMjC3CxbGjQhlXTtP5zrxNQRBwRkzxrcSSWq99bohKNfsHdUoxn
xq6B3HErlpL8jM0tDcMWJKcv7j13SkiQ6e/GPTatNIVNxe/pGVJQ35mRQmRPBmXUWJQAugyaGKCN
YJ7GIr7PJFR3/d75SsT4NcbCCXksooHnqubzKccClQNSuIMVlRif/1+BLHj+zY290Op5VkWY5aCi
FFN9nUyPKqKTESZe59bP1RMYtkjDE/QyUAkEYEDRpGcopK7Pk29Gm6RtEhrsAm6hFk2sG2o+xWNi
cPPq02pQEurYOelig3mquZmMDSRvXe3CcpM03SavfvfVX3xeZHUaei1Pgp0rxyeBsqt3tknaF8Qh
kaMd/iCSwhBlG2JAVscZ25VQz8QtDmeAtobSVqTCLsd0/3mwvZ7m54k4pT28ge8WApaYEImSWOXO
kyedQ6j2sfTqxXsP2iN+n/sibkOAz/efQQ+Wpa8MuuQcMn774WvCvYM3O8Vm1VJvfHmLJQF1zE7s
gKpP+UTFazWSKi7e9JE9m9wuMJ3GKmt5zCmK7cdd6LbTopPIgTB5cPrqA41/n1Obzsh3MwQroT1C
rz/j3a79V3Re5r3OanUMZcolqVJvfYmyB7pQwJg2aOkZrXwh1i1PZFskV7Ds5Orc0E+kB33DyQEH
1oP3xfQA3Va4cm5EvIwQb3NuZnfiNGXKcqSDWH6gZK9sU6G0A5SP4UpXltmaLPlFND5WHBQdT6Pi
PbLk0qlwnDBGIs4BJTUCylz4I78Iichh/OqEBZPPUStzzo0tSbp/pB3CKJoPS1mRe2XqDs/XeFbI
viIB6qzhGSL1BEnlYhntFfh5UekiETP9kwknRgFqfxSkZ26fRwGu8EB++ZRxiJJVXmkZbJ0OYgRX
6oPOQhE+rnfw0e2Kpm0Xc/0TM4vvBPkZJDxRXiB6LXuTNdcM+LucuQArA8LtDY6QLgos66Cx4sE6
+VT7YMKAGG0Xq8QWLcA/4Il/yGpfyn7cccoz1/w8b5JNmsGxuCgwTIMGqMfuN+VlgvziOe9gUL2F
v6l2AfDkIPD0oNg1TftmoEBiDS/5VHdKcaSBqu8fObXiVlTC+OdO6GIxvYASE+EKEvsCghW1akKL
6yAkhKD67dhp/d/7vKPCANlPf1FR2cIRr19RDNELmtN7+54bWe01EMUbYWggBZxc9aALnVdsJDtY
47pd+gUPUa9/5Di+QzMrc9EIftzCl9qrnzMyoBp0TSp1ZsdJCH9xmoZ0aCKs1Zjq9k/xR+961TH+
cV42nmvZUvgRz8knVf3r5IXt0/7+xFFoyNrHuRw0DWO1pZAwZg+U5+HN//PaU4Julg8hVGHvKcml
9rEDidyBd0VFuHJ1Z+DqBZ6GVPbCDcCGnxrfqqFE0XqMPdejzkeTBN5gYq/6eqiMV/dxwRjSTYLj
skDghe5TBeNb4q1YLwB11ooyJsTo5nQGr7Yv5/SVsljfL9QxTRhoneBFiiYSlc31WWZ0GxAzswKT
1GIO8kz/mlOBEiMeG5tkxIGXJ6MqH6YSFjkfR7zWdDuZxPvKsvVNKX9vqqyTCXu77JAhJ9EaPEqN
ifYa6+BTgP21jfuzGB15USodmD2QNP0Bv7aHFwLdU1E4yi3XKppbS/VROxzmWoHMAZgMupY2AlP5
Zv8SA/J2LckdzDlBV+/St076Ot72RL9SvWLdzrweVpGG64W7AGJQUcz5AB94/wknHOzEsMGLbh3d
FHEpV4tDvfxev8vqdkFyWND1B2ZN5FTO9pVQxTEOezxqZ9ePHW+MXRUg8Tp6WCGe2RQlXi7EL5TY
P/vLi3aaT/OKY9551+2OfUbW1PpbGX561Aquh4c2OC0R957TGhOgW08WRZIPqCn5Fhpcs5Ufh2Yl
je3pLqVsRZA0S9sh4B8zC07yITGTW8y+66viLPIYVQ+DHO2LR9iqURE4RDwrfsJsamd4Wo0uvyt1
u4AlyNiP6RwZvHBC735AtIDpHEYN5ULcl9jBo1FGvoHav8VCi2IbJsGQL/MhqbZWM6fU7gAdAIF4
opliFGuKORkwvoMyo3SykmoT8f4DOkZOJKcmiyn8v3mlPCAQE6N+9SCS7uahx9LwfNAvwDV7pnJd
lrUYrzAvVZAals38XQIjXwKSSkJio0uL3egwdNlYepBmdTmjbuU8bqlrnddKi/XfwyHgX/M6nlWH
kxfx2QK97voAZWpyiBKG82sC/3JPzD+OaLdlRUVUIz07LmRQzV3yXT2XnJl1f5k8p4rKQZqJz1fU
Jq17sMWk+towacj7H/6RqvCVqFaLRxX0wPXhbI6lfKRGNzGYthPkJHgBfDCisGEMjll2ugkljw9m
gqqpj3vPidNl157ozKo19rkjSWzBiFQ6uhW2acopLTO4CyTFIV9JUYhF9ukSPp3EXvTSA6Y+7Vg+
xdhAK+xrI3Tl2cb1FOyveJ6GGA/vCryNUWgadhLgQozZUnvHEYdzuBQ3QIc687NBssWFCvzcTqUg
lVWYKgX9STlCTGPLzsyt/BuJ38J9rJH5fT0rdPD4L6ZQGEQoKdJvWK3CQ24+vrtiQ81ETT/xNI5Q
jJpq8HU+yb0+xzs4rEDJsl0YYPDDu7ugaLLi163r6Cb41hWB3qV5Km5GfwzHiPuRq0kXsGcDDy4W
vlHwIlPbJwbB0NndajBu9L/II8UsTV3tG7Tb3jTGcGlJf3HmGfJtRmnvb5Ssxl7ra0PHB4+HRQfd
8aUpcGy1z1CFhyHFxQKN9+ZvMp6FP4e+h3uhTZiyPaNDA4xRywDcigwIY209A3fAQXBNHFFZEjRT
JoFD7lCbLGOXhWY+q2sfUptnsYwTNktQapWq0RfcCl3yH/Pezr51YkzsVYIH265v2ThEkRj+/KJt
KiRSnb99vsCTZK5UZ20OrLpVWsv1KNJgHdj0HIpSO5RBTfcFOBau7MXtQW5qFMjUgFu/73MGQPQk
swnBn2qNcNOjNGAHkSvM59NWWBCtkhtUdongKAKfQhvwJP80UWSPfRTB1mg091uUxLgosrX3o7Xr
fmTwLn0wK5nERd5VOsixoIh/p8zPkdQ9kqZJOcPeaPUzFAwzD4AkJNBdIloCnMRijhWswW8FBSWZ
/SpLs0VeEaTdrNUrAeM1MuDw6IHnH0CuSm/rAdI5NK8mAyhmnTzu7KwSbf2zQ7OpsMvNjRjXbHPc
rOTlX3cMu0oJMZp72H9XwX8mhfq/ENhBbyr9GtxdtxGJ6wV8k5CIe5k0zl35Q+nPfkfD78FnhFBL
4iK1yymQlL6pWD4Pebtj5jFCX9fhtj3/z56JUk9gVdPpabUS/wAyG+4ZD+N0TPE0buppLwzn7b2A
iBxu72dV/rfI2oZU5XR9i9Jr82Vvr8x1UOCXs2D7EsPVtOa1ga6NOjg4VKEj+DnajzluisG+5qkK
hhhp9Evno16XFxyd4nsMX2bM63UyV2yv9JmYyKViqTQbUrPyUEQZ0jocsF9e073vEidf6pkgyUAR
37Fs/ZqVowgE8e8qZlISuZYIR1cdg5Cjild9zLP77nyrdiS0uTT5hsQfdDdnVCVwQaANyqc8wvOo
b4CUSS+FTG75rsAoBMOGDe3y5PbPrTMbU1I9kOVHHFFi2BqwE/pQuXaHQ8YJV6GY8gwExnRi89DT
IdbsXq12SAuhMkqgHK5CuYGtRwZgsYRV1l93SvrVrgmeoCkgTWGFaRndVAyjlbq1LNYddDniH/g1
4Y8mRiIVyceehSo/pYsNlKWawABrcDqmuekOj0W9Jb7XYJDU33nEpPQ5uvvM/Ex/foMEbPmWm8KM
iOzrhDTSjIVJNx9yPseeabLMZlyPcuCq6tsXoFUTS3lrK5QH0HfKikoE9CFHG1fe55mhj5fb/2CQ
2TVqi7xMdixPQSCl+JHgIUTvnpkv6MBnn0a9cET4AcqMISPdvDmfPJD5f9QX4dugz8OMj8TQHHNz
stuPQYI0hvsW+o19Y1oc1R63W/tC2QPsc6ZsevH8g2Mf/jXuS5pXhKMdspDNIcINoCYA4GbDcftX
ad5lrSd8d+9aIA5VZASvrqyABrpiUs6/FLFNYCIVniHQTbtGShHh5ZChzIaeXT5CRhKt3rTcksbo
dJp1l7+MBDi6IZeQfJXxmqiZLoCLkORVfBWUxXxm3+MBeligPa5WyHaBHqUhzh+BrnQOgTuS8RdM
wMdGRYuRmNJ3qi6QkpP1pKewShDSXfUq+fb9kF5POHuLPPcSt28IKR5RgkR9UGG0tzPe08I/kMPr
T3LuBDbkAhA2uplyxvSV4aLrzYLQ6FjtMNHeYP0GgUnpK1bF5GSk6Xw7MmK+dqloVBf/auRlAaWG
WgoOtYUQpxpgKYRkehKil39KSIiAljCq+rByeIPmlusxS9DifIFu8I69frIfIolkTiaPkZdNFHID
cQh2djKVSi+Nx05bPGP9Kiirv3fjPiT7L9cS6p77wm9X5awgtV7dq4wZJUHFFYsrCeg9HlHOU14x
N0ZfKBBYLvhJYqS5bzOpuYkSHptK++wWYkBEVHxnQFl4f+d5wg5+SWc2EFCxzpBc5Mjl7PLKzNnJ
Zasn8r/6Zm03IYiX5kp+6IK3w6AxDQFQsev55QgF6GDBtjuBE9wT4BaJWfYdVLflUlo2ZqWT+b3s
OOAqYcHi3Xqz0ColzFIC8uX2aVG0qI0V9c3Tj+YywrLX7r4X3NAz238CQ3syn1+V/QmcjdxR5K+U
XuKFPQ7CCVRfz3vA7aPFxfGwI34hSwfYR3ksGcEVOlrEUbts9SHMjGKyv3MMrGpH9k7LPoEdsqrG
aw2m5d6FbCvvpBEApcLSpw8J0EFCs7PUYiodpeU6udll3Q0hZPvj1Jlow1rjdZp/tz9xFTeMIYd7
Fba33LUe1tfap9JlV0e9VlF1T/kR+5ZbOdrGmM7M721ijOkn3r4vMdsasqzivJMJMQ3qZe6q+sbi
RKT8yKfURRFWUnm7w2515IAl+Ynx6K2EEXQuES521uXDRr3LzX9pyTo1dVCKgjNYlXdvLm2kewDe
qUzwC0hsdWDip3PaK+UJD9mrxQEqMAf5d9WEiuCztdrWntC6JXf0vBHrHJgHBskWoeiiNW1+Sjqc
yKfby7gjrPfpfLk6rbW884xi8yrhjJrfBqyppwLIRHx5kaBRkfjLwHA6LIWex5MLHU6Bv7M6YOQM
HLf51RN6sQvQ3MZMWTc932U211RNb3wrDZM1zvYXmKNjqpHyyuNYHSFqEdZUcjHS2wdX7vRZ0pkJ
htil2QXatXKPBwmw69EHJC30yov5pdypdrQ7nmGDmmhu8ZOEZyjsTmzjgxdTK++mavwWVvzan4cQ
2eraXHk22pm7PMhpARKhRsfJSBpKgDLF0IG0sN7PVxpOxYwoZSB2VwdRScmXVJKRaKcJYBjINtny
tVmaId0F+g/ZwPWEsBIqFcFvgqsis+9NCa5CXh53LWI4ZzRgz69i6ptODgoe5cCL/Qz1ElHx8gNQ
ejM8Ns9mc2Dgy7o9qYMmcjkppcS+6IH95LQJb6YqWjnVrhAYpCGPYMNBLw1vbha2rt55be+jZIqo
uvcxm1w91Xfqs3IFll55YobQaWmSwoHpub9YoKT1+GY1W6IHgtKuBwDNb8bU1OBMr7v1xpJg9EYZ
Yo31ZLgmmee3YxbGT+3z2arzcVxCsD5tk92U5Cbjrttf3Li/qssiBRXY4/RW9mMPu9Itj6UgE7mb
CBiBc9GbBnYEyP1uI6c+LncIaI3lunUsSkPiHnlUBpRn1Uzykjqy35Uc2LCpU6GLDZhAjUqgneTI
ycmu7OX0F7hqgUfgR3qLs+8lL7x9HGUhg31daZdByKn2c+Eg5KcGTCVmwxVPtitWhmvrcXQV7Ugv
hwWyQSdMhAG5liTlUAM3mG9er1IgH2YElCQZNPE+mkIb7jRQaR5JYBlnRq53u2HNiQllCHjJyL3V
1JxvvAT4lU1x24shtfTHO+/ap2CVm2WX+aFYd/rpYSUSYqV/LyIaBcecAcoCP2U51yYWa428GElz
HZsFVwxL2752lnUpsNO8+/hyuAkRVQwN/5e9mfY44XbEIEeJsegsrRITDmIiYovaq5VAGIXgzFIC
iXyCZZKxKcjCEo4hv7iVcVEoCzAZFbO2S1kc1v6BTyD2oQ3C7RO4hHCoGsJ088lAV4uTaZthNBrq
e69Jz6TRYpwWdYFWirg/mOzqtdSSP9YczyFVkhjF8Qm/9DJPGgxzH0uGhF1qBWbjEeubRKUuqfXA
Hop4QOG9+Pb+63dH+mKpObuGSuHMPKkHUANEgsLEDoO5+hIWmALiTWJ31xtYU3yey8l3qNRtvsR8
sSBXHu4wJ9AjvrZj9FF6SQKS4+V2iFjThM69pKbDimUsrvtm2RUosO/bPoamE4s51gh8p1xCwHL1
2oM721dYdS9mSs0Xk8uE3ZIe4ESmRK5WddLXwGkGHuZgJwwxhOBfJDaZG+ldNJnkXIEHYvFn7ZKY
43J/FD5NjMg9F0ruFsDoq3QTzjbhjULf6D8B1KRMyLy/FLwnpM00ZqaJrlsH4MKbOkJSusS2y/Lu
5NzoYgA59SWlmfxssqZt1nD+tkO7EYZJd1/jcSxLJH5x6nQUBPJ7hcXtHFTU+cAhYQjguu/EfX+L
ZIEV5qpRYY9HFu+t/Fum/NkDBJ5dYBmcv/Jw+7+uD8YDLXXCEkvNykJvcLVkut8q9Y2CBBX5lKux
ZKtiyULOrGEiKjlix7Bzg05VC6gn4eAPBR6t9N+buBC8xtJx0Gk8G4OK6uDJq2y1eiFDXaCwRZH0
QWDKrDbmAik5Dzs0kLHzHgxgP8Eu8bWusD7vXv9J/uLBLaYMOJvLtAFw2rKKYG67trUyw9IByXFp
xyE+Jd5aMfSnf8d53m19GNxvNwr4/8qWTNt5R3OfWimYniz8M7r1pLJDKPbI/9j44iUL9UGouer/
JqlaVtM1vHEjWjY91JA7mVMPQmDHmlNvnun+Ljl+2R4dESI/GctkodEAoCpGmP/i/Nfg4rsH5AWj
egEOijsrz6OV7dedXg+zEkLmYVxD7lCLu9BD8RE4YU2pS8MWBFyF72UTzKE7yFwV059BsGuczQ0X
zUBs44cepq9D36aO4UEXa2Dsb0IiuGoGCNfzbp1bLGSeCc9lmOpwOKI4ujGftXqYWrZxN0JxEtR0
FbHboaXyjYMtE4UtsbNTzKdLHVQ6m0s/rMD6iQe3jIcW+cKYHFdypu4lbdQr9SmFJmNtQbCTOlcV
TMduP9xww8NgOu6vDQHM80jyd+5ccKJLSHhJE5528qN3OgRmLc3qk16LrSoCcKTHmQM7G//ZeCaH
Av5b06vvsLDLFok1FcE6IcwBWwxcENPbeBzepshgiQgusz+QAaIIF+5NuceMIsGWDe6C1ZzJ5Jjj
4qO0n0WKER5w/ev5jdgIG5I74l+z8F4t0t6epyEP6UGdo6BqGjfnI5ygfnH65Dr05GEE/VdckgSt
aTHtZCMhhJlcYFBKLQoZLotGV5fSLoNYnc6C78vf7RTr6TU9d9X5hNVSK8MpNzoIMnJh75VUeg4u
Y98HlhCNh8jTcj/doOwNYuexG9Obk4Y8f7HSj442D7HJbRF97i39mzxjVm9VEMKamKy5BiD2zc0k
vvSh/j2Hn4Cvwem04FIVyMjhUfPayitFp0E4pdz/WRcT2VgP9lZM1TsjuhRUGvaDhJhqOQJIDKoO
mHk00W93GKT/XvfAFNo5MAUMBwzHXp97mORIs8PKR1HmKiBWFvjsCm31HBwji3BWZdBxyUVQxRJo
sFc0EjR5uJEVPgQ+G+XP2B84AnYZzykf+8Pz3B7JIBlLtoLpHf/eVmKMb4EQJ+pQDCfprMCRjAaT
eWtNFXX1MOynjmRSlr3Nb6JXS1RLFfUmDDiLS1uUTOTi6GpIxIcBTgnpP/J3bay5Bchk/1dioXN/
2tbsdAyrbZ6fNhw7ZFvdqNTekyko0CuQri+T5S0YG4kIcX9vsF/GJzUfAG2Wtp2VFRLpmPqmZolC
vqdb35u5swF00SOshKI9KEQCk3RcirIw75CWYIcvszF81VEr3ohHJOI7RAAZoWRGuQhB0dCJn5Xe
P0r5HtbsV1WnF/aSUlIEUh3uTj6Qnv+5vzmqVSJE+BnzJRIrFzHP3g+PQ1jPCoTsJCBNQzsEqDXj
IaodPQwkYt34HWlpIzQ3VBUqEI7oILdnyX/fyLt5nEJmR0HU8B28345y5DozRSTTxCGQhnN7yEGl
TNulduSA/FtkkY3oSazKPxb+wm4OLxki0hmUC6Fa1IbeCNHR3Ed2JfNu2HQpWv6FE3r5yoWTVAFP
3wNFS50rn5AmeHvQ3BqBi6aYO5iwvwpfAWVjUu/OVNZ1uKtxkIurwoFSrylo2ebe2ex7LfuAxQC6
qDmmb4j3shDxyKJ5uXd2BpFU+BtdIoNSjHvLH5Gd6/6s9SeGKZv6bDhNthrz0ZaTwLF7o1UyrLmy
uzhXJLLVGHqF+Su/lKgcEZbN2g9SgXg80dtU89W4GnfSwdwh6s7GgCvrGAsMnNCiVh49b0RGrD0d
qsmHOKSIGMokhfs1CUXllz/NqVGkbQF6McpT6bfD3Uj9mZuwPZdG8YHgmlyngpmdg05W5P8xUgZP
iuWzj4Fa9fEeI3M2L3J9sq6tw3ip+8RDNwWbGhgSPj48GDstTKds3sGaBa0d6aWG6KyD892gLCE0
qOjtfoP3zn6E59jXd7xiOYbA8klJrFkRo2Cwk3UPUcFFb2mFjhZjoEJYbASOJp/LhnV6y3HFEP5h
RxmjR2/zl3A1SSPcKY5KU/BwDUPOkRE0nuAytYlxjp/JCe1gxC6UU/ZTvpe8E6DBK9q6Xm1BwYFM
Yt+5pcwkYGag1siTOvtAKw8b1Vn3OhKO+6W2/6OuTldFtzjdniRQAqecjGq62wkYX3EsnYNDxUa9
pdIYvUYPs0TEE5n+IhBAKYJHmdaMywaLpyP/8t/2WggBWLAt+v4lQjNqLZQIYa2EJVHumL0q9Evs
Wd5mKpQK2mTT0JB8e3i1hQ/ks1M/5Ybs/onizChF0ib8d0eZSbvLRcsZWEqvaDzenbTEHCOqyzA7
NhxEuFmWbHjLgD3F6y4uKJ7lTjtTOAWX/QcSGLUXJb1uPsAaNvlyR6yWiaIb2wyvDBBbPbPduk8n
0OrWMl7uy6PM1ZQ46durvgALgzM31gFkwBoBmDCu2igEaq74nnmY0v1XBz8vvOfHM9ojuoMPQUcW
WNmd59fX/hk+osO4fOPW4/sfWJ9xb3Uq1EAfL9UmKjRoiOyUxW0V4ThFBqoZ3AgSRZOGKQIRQu+O
h2XxwB4NbYCPKIbvcnKch1jYK1DbdmL1bjW+mGon0wQKRILBN3iwafxGb492jvg+fi5Bc0AV+Boo
srb8395X2JcFtw1a7tbWRgRGwPrdJJANvCnf803e7GkxqUt1eqR5BF62cKm1uMQUXqUvNOAfBF2H
W9nyfgaVbHZuLaFk/xwKcahuRp+QgVfApSbcWEQj+oG05d1Oslis5UuRGf9DN4cFA/nZSKpMnbaO
0ei5wvLVgIh5lxaQGbii+pA2G6Fc8AHnWC2z9GO9kV5hq2KkEr9gdv2+c7ZxJAylY0iVd4Ng3O0M
7ufLLRGapw2rRd1v7jlsoGXqTjm+5+YhgePqB0Lgn5VSDjmC3IWn8m+uJZ+CEuVQHf3RIYTZz6Ms
Luh30t+HbksFvWXBweOoshrpOQ3dQ4YFlmUUEFAibSTVEaeFU6tmAFjMABsEn8NE4BzuLr/BeQDi
lD6zH/cfJ7FqP1zFyMjPsjcXvN54KTNojxMvyS4cwycttq8PoQ9k59VAorrlTztjgixsX0y592of
W4rLhIvtRsh9hJ7vzN+VLJai7lJ17tyxG+F5Tj4AylZVmvS/VCtIVGgMQRTygkHVSxia02O+3U57
4PaJPqqwa4/4FSMx4HahvBJsNhdw6Zwk+tCXDoos/rdi5d8L/Iy62+dsC8Rzi1P8FXbW4ab/bKTo
MRS9FNgnHIMrl2oUiH62/wHwZam9s8c2ET0fuS75pXDUY11eezdXMJ3Re45mysdyWzj392xxB8mR
tvGtAt71zjNRTrYLxlr+fwjx/XUQKij7uAwG/kMo2g5ZEsDcVQO3m24Jq1eU4zInI2k+TIhrbUTi
m92oiF8+bQCpThXzPZ9v6E7EA8aXCLY5of/ZdmJmr40URkZXGjrf5ZwF4AiWZRck/NwxruPGxp1n
IxospEn9NHS9fZEnZpVzxB6HJYPOAPinUA49DwMraWHq7ScxjIgykzCx4vVggT6rYJ40Tgc5AQSl
MzdorayqEs8H432gUDFvnj/zHBZzXzgAXsUHNuHYN1UKXLBpdqxJAoWZoJ/J0e5MkalUes6pX0tV
5TT5DZlLJ2SL+F9oJpm3V/ZWdkaF4oxhI/d+f+Z5WcZagu56NSD+HdAPkGPanOFMS2QaccEr6wqY
tYlQCaLyuZnavdaOzO/WMQa/IcqnWr8lipIyAxyecTrz1jWXWyPHCLJx3jotX4zNmFaXHKgWTc8r
OeDeoviejt3qFt+9/4yTNtLGh8dnYkBY1IjN3S/K8kWdOM5lTcqCLQbDnekicsXZFJmHG+GW/IP7
WNGLsujlFOfu1RNcG0wjeBnUyuyfDi8kZlWP6OBeKMoixZI7eCwSWbS7+S6LtUlxrE3aKlEsBhV3
Wd6/l1wErQv14MT2o5o4NzTP9dJ+iGh9aLZxQ1hcYkSyGR74OLLwa0J+uZT27iYK/Yi4EazjRs2w
dnbFwiJt0BQ1IXIxzNYJGzpqOtgg5vfHxrWQmWoUzdgeRg8KFSdWTQ36JBYRzF5s8gcCkYOtZm1U
HAml6Bms2JSqxI7M1ATav/6aV/ecU6wixuxdCnqkW3OQof0J+00sd/NMlM02b/cYb38a5ktQxk8f
0wzsVkn7sbAvDte5P03ssBvv2oolTEbBt3LxR+QbSS4+tipIkL/ueBvjY5G7UK/o/nacpZxvuNKG
PR7OsvxW+4uC6YpRG9jyI8m+EhfmGhnASEDsmQJrLkIkLMgqc7++UGbq+wHDxNJmhQxSJS7zmxW9
S7LHlkwL4qd5D8Sk4kXNIvD3EIbTSxg3V/d3eKy3s0rryYZO4WNQetV44rU5uxZpAPbRO7FwGE/X
RLbYBwvACMacgZCrlhYnoce6JfUpaCFesxVrhPRz3721d433GTOoqpDc1m01biLb2hC+BfTjVJSY
ZX5+/iY0ecoy9/K3MiWNk57Iu6mfCMJOsoW2M3wtPRJR2T4DE3ID4S0VlhUOZJsX2CNZLWw4tPqC
iN05ZhQT62mTTz7T5QpXJxtcdVbwP3QbBC0H/09qgKlVR/sYj0Jx4mu4MLguQ7a7yS3jt19B63yD
Ym5AMxxLXYjHKXh5efITdwBf2LMCNcsnNCbctROkxBBKv1S2g0y6UqxrAQ2yemXRcNE1CpAy8iR4
qa2ZRWOBrWCx5HGm35gb+Nzu+amzx0mIdzpM1XFOAit0yExKaUxq84PPZYWORXGROUdqiS2K3mg5
EDUwLU+izXfR/v54Vhdr42vjnU6ltzqE3e26KgeOc7+xYM3yTDmxlrvIbKRf9ButuVMpj6blZe09
N0wmTK3nbHdbwf01yrquKwi1KWSDqX8flsKwozLe/uSzx6XnE73QWsW2hxH5W91AyhWTyfGueufK
clYiMHThcPu6OZyXZ8vDSWcYAuZUT9ZJRWCWL6oZillD3Oq0Iy7Ubvwvenu37zyg6T/FWenLoovg
H+EoWB3aukxhZlOac6KVx71mieyC2cqa6M+mFMWu/mibv32Rg8R16EISIyGQ2MgfFtA7CoENKQ/g
VnoHoyBYionjJHR5GG0JIyx8+K2vj7L/ed4hxP6TsvELLellb28n/I8RrTAAlGlByIhcZ7tzSq7f
u5iMKDJJt3idkly6+AKjyLsOy2kdGZd4dfqD+u8IiB63CGdImse4QgSk3Qne5aFZDPns6iiyAb6/
FwFJqjrF8KUBUudC8qtdDF/0+QYyL1LJBvmB9RbtSXHOJsoZ/vZlJfyX9ngKfedCYgmVvtGTtCAY
wn9eMT/j5mYJgh8rRi5v7IV5UrbEvVnaebUfuakK2nyZZj+V1Sr/0oRkAkl/yC51RE+9umTPBpbY
PCwOlxNDXRt7t0mI16HBid1Db1cqbnECvfacjNm02UaRDBt8UCUst3w8tcx3Btz0QAbGdGE8hJYg
fFnAE+nE72dqSXcj3/DrDcR8tLAcyseLY70kASfrp5hyyQnjf3odVSw918k52/JKGlIQivXrfUqL
whx8eTzKbvcizdPQVGkh7OskMS8xlQb8QfHQv4i5IgeiL3JqsfJkbaQVjpFaZtHecGq49AoAy3/T
YVpyHzKtqGY7JtaHkpuUPcnHibnISBCjT2DWuYXT8Oa3tXX4UPmbVppf0lhGw9DTPqlfU+7Rzars
GmGoYBNl+2A16pnFHtgRUber0C3sRXO7KqQ4h5AhDfkm5b2mug0WjeFNR7MJ2iHlNRAi5RGUL/Rh
KAU5yugdQp5J94d97LZFoAcdRuGiNuKjFyQ5aRbjngYNcOQyVIJuIourhTns/8S7qYkiqdC3FpC6
QzQN3xOhr5CfDjVdmWEkreTZtZqpVLsC+PjRJJjko6WgfGIz6udVGqi7Cq65bXWS0ma7aae+DSoa
C02aYq2rSeY9qDqWwiIndoqrpDqwJNc4BR6qUZyn6dcpgaUyfWhKJ6ypLjm6qgOyh7tWInRWNEKq
BxWgBIReVHfKS9ZXxF2MwfqPYgO166+fVPZWvmC9sjMAmwFNvFfKaVJ3bU4VtPk6p2feB2HCcUQa
AHEc1aIpW1w8FD/lKTZIhbSlj3jA0H5+FIfCU2bDqlpt/OxEOJ36oLaG0zizspwGFWW/SeE3jvQN
kZe/Ah6S9t7cth/hMb3HcZA7NWTAIJQnKbBpDCMnZUIg7yvdKQK2j8e6BMOacDVVTFfFZvxim0cV
J3HbufHRjvzmFBHqnv1DoUKU3E1sCsAS6U/j22Q09fgZUpvuRJNA/vGAKanI9nnJagnzRRVO5ukn
bciOa0hIx7+CdZ6/VU8ZCB99vWqBDRkOQZ59XpMOOrNVesqP4KhGYNveINPAxAJE1isYADMgCSQO
HOa8ZIoY7/Kf2NCdhd6TIysLDtiWsaJWj0ViIM2+aQChmUMYo4qaNlni40QbhaG1YLJtKYi8+WDd
7usljiOYDt0EX/Vbaz5gwsnAeoJqwp8vIwGHNBKawgaPow23Iqg6nyIT6gnAgv1wJ181LybJetJ8
h7rgh1LrxcCgAWe3VNYjALfaYV6zEgrKyvDyKO/dBWl3H7+7JLbLU52ynsZvYwc38HB+tL8MvvNS
+8//aa0+3XM06ZgA6zecTqj53+AZN1NmpdRrXvjfPLeIvgb9sV9GLQurW5VvjbKS3r+osC6SqY4o
ge4dmjKIyKCg2lcGkynfHlrv+pyJKRJ+tACTLIGZ/wqjqb5VrbWC2qsGSJap+HxJNME+IYTkwVka
ksgmKF7NQGyhrSPl8PznaEpMTbcFudQbXVtWwj2YYqAi/7gADTyZ7CkBwnSYUpTKzGV2nYKDyqxP
5ag9etLmZglPONOO5Yyr7ObTYc7S7ZXQ3pzaWGgZ+acGsLfkLcAsoFDofR+DUlAIvYZ6iq9vpO4j
/d0vZXXn9LBtkaIWhT37J2IS/yGbWEa/Nknx3FCPm2DrUBigEO2Y8w+F8mABzhH/8L7FgaBgetUM
gtrvbDyJji4EalMy1ZEESVev64k4kBhIV1adPLClO7RhBoAvuZjcmA9Ctl2Qv1STXsRBw35ZCu0w
chXeHgXFQkaLpyzI+BAV5qDoRsGOPEWOlLwtxpNRXDm54/Lfsyz/TvzfLIAwP3cb6zweOtV/3Ple
BN0yIWMgBLL+3blvFn+DFjJF6ouS3JGRpBBCY3Q9a2FjgOfz+oWHDbt+Uk419PF10LVR1/ldSO2u
TJmpspfUGzjYk6wW6rzbYg5lPjSudgfHzBbrBTMwxu/ArMz8+cTpJS3l4eaDDtpRXg4gxH5bWVCm
AEmSkf0tlYzNDxifMx8WEtJjqrbl/KHea73oTH2AAML8ERj6wXwiO0lQukLe6ic6S07X3XvaUeER
Dkf+zdMAp9wYFVNfjRHNkeW67+coxnPq1XCqW8DK/4/3j9dtG4meIvPyDHosI6lqfD14NWVwu5Ic
7hITCOU/Nn/HGYhuZxHYwVdcEORfm5TbMuzicZS3HeEU36q8WOl4ucw0QKB0dalfMuHvKaGLlZYj
3RXDNpmCmYms6DASc4wz9Wd1ZzPuz1Dhz0VUba4fAY31/nBlbbrMqb3QdVUzT2MQtKlo9ar/7ri7
SGD6COXHPmNaTC/iOaX96j1IEVvMzOx3heYNrwAxqL38v0WRcZx316a806D4eq64GBA7loG3HGIg
QfZQHFRkOZnqBoFwQeeiirJ7u9cHf8+Hj1R12ZKFBy/S4Atw+0pfsWwf4Cj0VKOB4PMHb1UWTbMy
OiMVJTbGN+z2e5gCX1VVm+1wwoLrYJtcmrFlv40cEgBD2KK8jrVIqYhDx/d4CdnWkEsRGzcAJfzY
DP7W0ri4bYZ2Cxsd0W/kJ1Y7oBJ6X/hkA8NJ5tpZw2JCCY7A8xqX+AMSn3md0xdgJiajSf1a+Vue
LaHvLbAWnMwdH3hYsRXDQXJXA6dPictej+/vAktP0PVeHzxs9LyFoZheBoqTL0rMtBpw5w2k+Trt
9AJAVFXw5yyuE0OUcc0Gfb3aRStI/8vcFNSVgDOPnSfqbuvUsTJf/S1skDqgiolF2aUSxS945Nrp
mTcp12rfgig7nGsn8AhBemgbEcOrCpk0186eKbghhTFA4u3aO3UTNEcTKVoew6hqhp+K1HrT8iWH
MvBtzZTLVfQ+iHwQaNRXzqxuW3AYZLzK4126vkKKuIuc8OM+dgjo3Ia+yl6jsGQKqWsXXGwdLiTY
1z5DPwmYH8318+d11zBWZ6Hi6nwEVuuwzcF4sBrfIUklJ2XTI+zl3F/6ePP0x/yFrBamW7sx0CyK
TEYBFouBtDZ4e5Hwyymu9M645PY0MuQzUznwk4LysTo6m0bkh745ILwLHmoJxum3kTn89wbYmE1v
QuKBIabkDYLEhHZnjRhhCsKIeZ2V+XyZGmCkrdNukRRxQazC19+9MZYQ+lIArwckXSIHlVrAY/KJ
ZEPSMlCj42V/n2rUtyclfScgYpGvL5WwshBDNpNYFU3QSIKSMf/Rtlu4ptCL2N1flPHZHE321P+x
AhLlKyap5baaQbPo2HXesBqdtBVlX3WI99+67ELr5L3wkG/8VAqzNhfUR94SFE5fk19ZU4MmL4sY
OKBjOUwNur0gcHueFzRWnZ+3yq4cZmvkGz06Rn+7TgnTbmmDQGfk5n16KkIrxxXRs/8zmsWMq4EW
q5D3UwVe3KPp+tlMmdpJ3DK/6HAP8HZ2AHRMHAWC2f5uesBl9TAPT+Uk6kEF4NscI38MnBrI32xK
F8CEDT6zXEloV5np0yx5ckP6jIBqNH7zdU/So6sAVsTSwcjQGmplnMyfd9M/8o3iL7cbGMdaU/3s
fYG+8Fwp+S7UjJQ7nEH245ovhtAwdesouqK+cC/FK4IpSajV+LzXFpG3d1/oU81vjacWQr+l2KYx
B5f9Wtqc6/nWo2aSyJRPKt8VLPI/SGXC8NsScrQ5dTUYbjSNYVifVSF24g7rDR2UN36Kg1JvP/vD
UbefhAb+2Om6p1KdY9dhnWykqvi6qIeKYRffPXVPV773dZ75e+Hiz6XmxcOf4XehO4F04RwA2QYh
AlB7HqNAlkA6zYb9RcqZzQ69MEVmc9lxUmIgL0MvgU2dOObCWB7dzEqZ/g22Mq+z2g+kh20whzGB
CFwD/ub2L3ik8IkhUPaJ840VV5bDylnBgX2bkVecZPF3O1LuRuy0chd50l9/MdKraSHLHA2P2qM4
UupwUt6bP90a04RaBFViFtNSHHu+KVBefuh1ZginkG2JSsdpwYwmMR3dhp1GvKIjgYoaHUo6RIKw
1KST9nm9VJaTHyvW7caotoLExeT5A9TSAHBCc9EFMFjLABsmdBVP8+Nq/xPcKSP0VJE2tsNUEmx7
VVTsxIXk3DE097LCeKIC9Rd4RwVhg5c/gzwPFSPMPSB7fq5tGqm6x3VAg0O6vRx90PvbtGR/DECG
Y6lt7WmvDnNQQ19+vJbuyrZpNh3/uMpJ+ftfbV3+RygAHWO8QMHcW9XibTc6tHOLwdl6daYjxQoQ
ISDrcPr1OeUTWafGfOtOgBK1UV3AvtdZj4GZxQFB2RWNrgfff2Fmjl7bAQGjkkTMEps5ZTg4gB0w
mQDRCcx0cEOKCn1NEhrC/wEmJwC61jIGxQEy3doQAXIcHb7bk8oFd5RiCgqycMQT8KEGiAUcFW51
OvSWyeYEYh407oG9uGI4Dlud++9natB7slZceBR1wt/VF2UaPq+i0iulkpMid2qbRiUsJH8wgnws
qyMqdyQIAqstN1hiV/wbREBb01oJoelx9sysJlU2CM5z5ODByUFNgOIMMWl6jDWPEUI5JDG49jHx
rxEhUDVNnszqHlUgupymIFxJreaXmH7h6ypLBccW+Kxt2zgAMKa2bz9VGn2NSd69sPNTdXpQCIYR
5I+2TZkQpPOznjwpbZY2h/gN7PgbD27ByPL0r1ZMdblW04dTpckQSpXXFFkNZgZTJHxUuFpqTSAL
2eBkRtErLVPMM9e4//cgbZYLPOpHt6WIDVcJx3UE370uFoEE1DJzV/VlpF4w8Es7/U8qgJnBPcPI
NACV26ROm6I8HuTRwfQXLEZxC1W+gQGCQklV1p+s+COk1zIMuRcqDcnLx+SAXy0/t8zpApG2uFd2
JvgGg8ZlnkXsZWSRDAaWrnRQ+2IqsmgpwKs9aWpAfFJLZnVVx5X6ApVu6xfko5gqmQr6VeRTBSDH
/g9pOHD4s0gq9L9vPyD2nrxKA8tbCwRUXiZq9UwY4SHiwgkdZ/MdkrZFHIyzoVikL8N1QH9J1D7u
XE26lcMt127s/kX2KJw0l9w7U8QiSuIYFmGciXw8g9vQUGR8tl9f8QPaiX7/K0BykVKyeS4T/K0p
R3oUeKZGrmexcuWqtz2Nm1g2Thx0uxhGM6kfZ4qmxj0Z5KEDY9tsnExRn7FL6x6Daxs9wEFj6gFP
8Jyj1AO/+8uN2nabJfYo1PaBhBMfhgr3N9VYaT34t3Q9HFcnJs2QZIWmr4owW71984uqlpB6UIJa
sKcdFUVMmMD5xNBn3Gb1jct9n2B7S5FCexFKYKm5+GwtXbCVF6yzOco50xX0V4dbFN3NE6Hauzsx
QaG0VQTLVMR1tcUjgqVWqwWvl77PD2Kye6kkt/DgfTLJVMHU5qiO3NtM/11NG2vRbAVlE66FtFjp
TEjbJ6yfcO+AYNeAHB92XCd4zwJZOmjWlPCkPAv0mtHozLulfy0wRX5FGmAnWkBQbyq0gMsMLGro
uniMEqyGcpOL0HihZR+HlCDpxAKkg9L+imiSKodxLO036pdbUAAIfwe7yyPSK2aHQYb42HbIiHyR
4BD1/qYRN2kruYbCF+gRZgNCjYY5q4jTd2UrwL+6cVklcCfVQ/0Y6eBYXhbe2C8gicfuqKZV2FhU
M2GQ9p7m/3FT3P9AfFTf7wHaFP2xBC3ZzSCwQkxBf3ytW0+vuaCSGgHVLnZASQBvD2HgIf2qzmT1
mTEVaU+Y8Ne09oPdm2T0C3u1zW8X8GmZhk1BQzEsban3ovPpmDLuBvLPkBqZRZDf0Cw7ASckh6wz
mAvX94No3EE586xoM224CS3ppM9ZSPcpakEQV6EhDLbvFqrZhfj/H+DqED+llxGUxlO+tbLToajF
7gjNO5h3V+JR8SqZgSbhqN2Rpoocew3OilmBrc0nnB6AS2wBlR4zAuV335dOVlucTEUvbFxZL4ap
MYZvOMnUd74w47IqfQ9INkZIF8YifJy8I0v3l2KpDOf/We/J9P/UYk5g2nlA0SglYogkBv3c3UXr
z+K3eZaK+z+Zwn9r+jVBd4NPHqAqGRW3/PXvZsFnQOCdQcgS887ptcgABc7Jq+etw9L1UfffXjJY
fa7s+5D0d5qLuN8xCsNPVdX20tBYYmEZ1VcPiSZUiLSuUSttkt4MQX24bketJbUN4V6KUR2c9P4O
4B+k3S0Bh/9BV+PL4q2S7ThOkwF3NA/zh51MZHx6TeAyZXmyshTIgfBoTBrq6pQRy7g2tin6vRGA
9vl41gIdvmqRNvq+b/ogG92jBnXVkzWrp09gcG4HTPWtKUXfr1UU6KsyAggpRUiuUPlqHOC089vc
u+K+c5tkJIJuUCfaY8Hht5zL6i59cDJF0nuMnRZyFIuICFGU+yGPDZ5MyS6GOK9PdABUVztsgCP8
gOxeiocxzE6AbAHoB8+jwiICBRzIMdWgg801CpdcvNabF9SkHOmG5j3O5GstK0lJRoFVnbhGPb9D
oUDABP/AU4M3eSs6IRWmfV12VmZi9vhEyhS8xQ0Hf/OZg1MBw74V/srV4lEJL7G2mNvXcoYrHJJP
zUs435RpcVLm2z+8ABic7P11rZGYQ4OdyyPQpxqeNhGMwKvMdSiuvmCtkwAuR5WW8GkD+9a++pNy
06NKhALxkNJLokGYjp1FyWdkWD0Y10O1oHexFBH/btPTZkkb/iFLZ3UgomoCAU7IXagPx7ARps+N
Xax5dvcKnWv7UatRJZsN1vGbig3BrzuwRzhiNFUN0N0KAodsaGnResaR7+LxsC6POx9LUM7SStn2
xz900W3i03K1SYaKMW7HkLU1gTprs9b6odWwMYMJcyYWxclBDAMFkx+HASkZC8q7r6hOeLobzBEs
/2Jt/XaR/W139LQpeXcRYZlViEZa+fIAppCeS+atmiveIZJOApY+zbxcVZkGl/FMchIDwNuJrrgw
L+EBdY5eSOdSmwiQAAcBG3LodEeHgV0IWlutwredclOvAzj/09zu12UPE3lTDzSfeu71lFPDAYUA
gs3poKLeTSwZOmjwfNSFbX4IzuMJ9e2FRLFd77z/ORWi2ur5n2SGyvIvwFLpdEofWQHfpU8O2cd/
vl8/4zOMXJochz3qZ5RXcP081KRk/ECag6XLi5J61hT0jpHwnwbusc+02aUbs3kCfudCGQ1gL7Vn
mQm5hcl5O23f05pcJoC/7aACYQzYU+1pxPzNLRSzkwt1eaThznzvVIRZQ1An4nsWRJN7jNdYHnFz
Q+7I0OE0/N9U1q6ZuC3Wtb7/Ys1AdJh4noYEOyZUDxTK6CP27jgtSrHOuJiQLorTidPV/2nwySBY
KN8s/3PS0iVMOFVh2+93C+ywKFpIlwbngQhtSj5U6SuQI+LUVmv1nUJEfxmOoFcTGIfd+lAyfcsj
DzBwg3nYq8DyCudMlIlP5j0Tfgp76Nm8EElmkBHsC+bHeJfc+hVZvDyadyHFEYU87XcscStv91qY
GEPDZZ4SLaQEyNvLLXWTfbdkLb6IgOyN6vFwRevoep/hTxoJqUAVCTV3EqLRsTjSKeakZQ8O/Rax
dE/PtdQE21st0YqgOODL0JM4yje+RMaaCjIqk+kLkVdxpGmdQdUZNaqEu+omLwxtRTIDDzUY3+V9
LFGuQ8s6cDFTBwK4xtJRdInrfx6Gjefr/rZDrd6kJHhXoSG535BB+G/MPUMskuNX4Uowc6FtKmeA
bSlOEc9dCaHRNPVQYMZQu/V5jt+nI0KviEENpKsw989DqcahmJD7mKDfN5AFDIEnXbzOUkTTnoV6
BX2a06TaIpC0JW/EeI9QO4VwgmlVPKze0Er9kKyeKGmNzQVaMNcl1mRO2bTHNrv5j/FHyqQina52
xGrz8+7WnUs9SVLfp2ZS4h4KMO77diyvrzBN9UTtTk4NadLr5DYv8bWY/2EG/9Ue6QZCEaoewyke
4qK3eOZ58cAWmTt5zTOYzVMP7QoHIRnsyeIYzVvMiuIDF6SxHCzFn1dAcsbDHhjSpPKPZUaU5nGg
7+c9Yz6wBKTT4WCK13msFYA9UYrSB0LJOBKD4c70YpE042TrCFuoFVP0kYXJUux79vqwDNilrcMU
9xzEadFjeew5RYPvsjOivks191pE9zYfh2aBpwvSKtdoTd8gGHzrym7N08jIq0oPt/RLtQLy5pMe
xsnYtOmCNd9a/f37G7qUpjewrL95xDK+Wa2I1wJWOqiBJN0HsxVtj77OE86vZu2uy5c5mUFKXbV+
srJqvqyqkYj0og/zt2ULA1IlG7a+8+UdvkUgjATjSEiA3iR/eHebmNE9qAbPVBICoKQtF6yL66ph
ryQFtda4tTQLjBqNdaGrQ6pq+JWQXX0YYdmqBjwPw6eF8OH+a+ODc32zUHGv/cZ0I1maT5BrqMSW
aJDfBau4BAaJW8gvJvNfcefI1IDMiuazlBE3bM/6/EZmVvRAAEP1EHV4Sw67EOFrrLFBEvT00ioI
ZjfC2XKAo/S7F5gQRG1iNpFj1GSiWd0v8GEW3WR2oYDxxtWAfcGfLyWDPK2qRoTm9jhb186hxCNQ
kls5XKZy34I2xSc3QRBGm1xVu8X6YrVraIAuFl2EOmtZXntM4Tu12Rp7ev9n6vYrtHbAMPUcBEF2
SZK7fmh+mxiXbljyoLlQx31tta0Gpd8AAXREiGx0aC6BxxCIjDvUayqOn6PcMHoFe5v9EFuXWdW/
6OinI1QTdsBpQpqa7kmH5jPB6WxmsuuKKlCmD2TR0cn+2OYhpLsaK1WBKML5JbajTwYUV8at8tcD
ERZ/i7CbtSLwxbPl9aNRkUVNpJ9cHpoCG2j/aOR7xkt3EfD7WQSmTOUZ+N0wPTYXfX2dtfW91dlQ
Amcv9GJSp7ldqZuVtDgpJkIuw4Zgit1BgF5Lt/4AGGYpsAj2FpHXtpaex5NfFzOAiCLgq6tGTybf
LSDA9KPXVvexZlGv+V/48dfZkj0xGG/AFhvvDvjG0PdgLj85WTVGe1k2bHHlLAWb5nM8gRGJc2Hg
RWrbOdQ+HDAtZbkJu4VT0aBk1Ciy1kunT1cgTOLWTkeNsSuY4vgP5nVSwrWF2bOHGG3a4Qenqidf
07ZHleLkUY8Y5mOJfY2iU+akrrUL5abtSuNJNQP8EtY8dAaHcjXttMS/AcmcZ/ph+e4vQ53o9xW4
zgVbm3njpMxzTB6nBgiLgk2/lxlwPGaWssWDvmtYBkTHI3og/5pZmpBAcnYPj52B0rbpFzMMaVjw
cemPe/R3ItcpPNl6VtWEsth74tkjYqC7TtXfPYsNagscWSCTS8QTmBrfPZeHMJd/f1IXak4lWr8M
ukpypOYVvsZ+T3kCv3tFQPiIYvtLeomjidUKPr5SovMpkBXKMxRdwdSwKn0liZYw744NT9wHWu5m
8/ATADtB7VVQluQnWkFW9MfNsbCjt9dNp1VqruVEG3Nl7dtW9x66XdcJshSugY3w0ZXXx4F1a7CP
YR5gBIgf/GybzZBsmG/D+hqhJh90+pYhqM1lTrVU66nfGU0zuvtoUdMBvKjrSXRHi6rsOTg+S+m3
wgIPDuo1nClpvRcA1ZwAx+4yQ+7wnH+41RD0TdVcobZXH9N8o5pwzshErHphtQgmTHbJJ+pZPJ8x
sEuW4iqyWXDOMuN9d8nCsuiNdM3aorS2928vfoL+i+zOgxWy2JjkfaDzLpI6qxetQT078mh+JG4O
8whnqo+cLops+0Cr23lJ/Ss93zjZw1g9L7FziT8SdzNnw9m0vahL4tqCiW2qF05oZzQFCSZYHVoA
E8QMf2bibrkOGi8Cl3xb5Tg5Yzc+ePtE9qVpkS7+SJkyB2HA4WcZJ6GjeAZK2DiShcGc20ADIkFC
wGerpyA2LSRwKGeFId+X9j6IEug/h+pxYbpuwX3IQUq3d1lNMDJ23KN1GfL8XRE6VU05Bjf75BXx
m2cWSXjZXFfvtfEX2gA0Rz6CbOYeYdBI+FQiZVP544kyGZS4MRBpuJJ9epq09kk0uUL9XqNYDqAt
B4kT1AI1nVta2/Gpwq7dmLSekj6B3qMjd1IQASjmTcbTCkqRHSkeAx6GqwreoAs8xo7gvp46TIO2
xx9vqh114w6KLkpBryPOwsmBb6Okj8MkiSRBx6oWmV9IgW2slRC/k1UEFrRA9qE1x2QIn9gaRtq0
+SlFnp4iwN91emNQUSEmJ1ukLsjyhRDpql4bjJqofwG93vkuudK6/Bq73E+ADN+FsFDcleQdwUnG
iqE+7fKIWq+PbzgPplWPM0X9jzn96MPgoSRG4QBfLuEFT/jf232P4Iwj5Rs0qFD6D1IkTOwXYVMZ
xRIzTMPf/XmtbXTTAkCVAQyOgYneFcK9m+fO6W42CjECI07Jr2HtstJBdOAQDc7vn3pIycg5wEFO
Hh9g6ol8iZdKqZ/ekOuLmDG0K1JK+V+zR4qoIsJyZHxZxeD1t+UBUZQVQPWQCC9y9qW7QJ7JZcQL
rggrYjX8LhEY/+LPN4t+lh8Cr7sxrZGsoPZVwFFsoSL5oFqEnXCOe9Z008lVqsgVPZqHC5f2yUnx
v0GfdFxePtetf5kSKmmVqJZ08C6nxpORL8+Eww6VeFktaIBgoAQZxQpAKTYo993EgGFytOnh2Ryj
kJj1PkaFXsShG91s+NV34h3MW/PEr+oyB003yHv3sYC8as0KsqCMTlgMcLyZvJVPsind30L0fuf8
Yn1HZKFW6i/HLJIp7YyleNb0sdy4DnS22A1XuewImAytjPsM8L505Ls/g9EM7HR6TYs4DruieskD
23TDog4RCMdhLQgNsZ7/WGcWWmZ2C0k9MayYSOBKYb55SBxY/+ytyqFkuiCqqS1OEMV4+Q3We1Hi
i/e39jrHXyri2LKaaiNoMt3m3E6U1Q9pMCRTQ5HQdr/2j8pCvcr0LarcSz6vewqEmd1R3n55585z
NZPyjVEuWmnrF2jmEv+riOhBXQnyLr+Q4vfBlRQsu99oVt/0VoUqAUqbcLXbjBToruTa6q9+FhwL
sYgUYWV/UqGUau7k/LU0XgYW9r62+Yzx+1p5BWJ/HOkEHVxUEvGeYjQ1RswmjqMWhw5Hw3jRqniA
8mTsq0uHrARwNXLZGVGRo1jKjqif7BZyBOQ35RWfMBfvQkh944G/F9DbosK0qw2fOSouARPo8HK9
akSCeGe2Y3YQ/E6r4hOrgf125JjXp/GqeiJse2xRMritt18bW1p415kFGGEu/eNyMJ8/NGa58E4U
tlZV/WLXJAnb3PF7bU3bT8cNQx9jhY2NDrG4RLyvh7c/FKV7ciHq8iPUjAv5AW8x/S2EmQGXfavm
Y7GaAL7U6ykicrVE4siAt3f3i9E1u4kjn2e0W/kp6Xz+bPnHUvfzNKHE1V/YqlZNQ8j8myKGS3V6
btbgHHbVArBf410qNfKMjhe8s61DECdoM7eEZTvX0UU1HB47c4KzbQOW2iq5k9jHWb01lJwL09y1
QEzPvbFpt1zF9Y9E30Q7JHlw4r5dk5jqnsNEXPXN38QRGWfWtV0PU6oIM9i8Cion+jaiv2q19aw1
IGtutSz6zIeOazG/gdyDgRPct+aElysdhPnicdLZCLZfY5tMEwZ9Tszp2WzcSkRbl9D44ImC+gGy
aNh+11l3jI8sgCIShLPu/kf5rYMc9OUyvfPJMdz8Sjah17CP5IsZWSkDtaRnAhY9cvnwvLoHXGA/
BVCMFoZ8EIvnXsVTlvw4Hb+p6PjREeOn2grWwl6MQ0qPGZoyQqLHqcSakwDcbZysyxpZe/HbT/Rx
BuABMdJJJa6ti3P2mA9wScvVSiDv9zzzuJXPI194aRn4ExpRzMzX2XIsarl6CX0ky+XO3EwNUnrW
qTxzytsTyolr5YQRkJSkSKfbKQcJxBLTmUisWX6M1gMbpb6AjuqFYrfTTv94NpTR7+RB3E66JP1g
lLrM/Lo7JdpMC3Z4kbLZPATq0VvTaNOGiuWLtLth03phiwhnyYCx2I0kYncA+9WKd+162pxr/M8n
BE3VhRrJC+TV+rmZECOXDbcCZ9wIs6N+4SRJxC/EoEZU7nlTaHERkbYf0EQ7z79QrgrsKTTekTkh
KPJ6gne3rvsw/X/5/sXpkCBVuzIBYBEjDc3j8UTm5UHkkHjBYCQJq6D7z8zbGekQ0vAFkCKSk1X/
DR+DGok8oP/p6bsYt+n8VCsRqOllkRPz/N6+5U76voRiSx6BK9KAvgIg8AgiZ1ICsPHsmOhDfgNx
Tet1btfhtX44zcnVIXwuqaq5YtAyvtpLGjGfeGvnrWyCEX0BQi7T148Y3KPEvjil4anaqaYhGgXY
WKeA55guEeWfJIDLJqs3mu4skoB/S4BRxzANfiIiKibg5tKcEfn7VXauBobZPzawN/rRYTAoy6we
yOZcSv+SdyFV5C757rPQ0R2b9km5eZ5thXOzq7QgYHA7wDik6F35vAVSSsrl9XbXFtW7YiWf2vUG
X62gah6Ddve5DxxJekRuBaFuMsRt43GOmvfSyKQEbmL3JAZK/FlB2bK0GL0szNfkxwi4q9A2hpeo
spuJEgS4p8fS0IDe6vvcs2k9SlOfTO57sNCyc4T0o/scWBEcOMuS+KdOwFDEsPufVd4oxwC+uPfE
vnaPK9dPoCqQvOVBQQ1CTc0KT00gaxu445N+sdck8ljmJ7p+/LZCdtyLOHq1MfFAZgcdMi98Tk/0
TkOOYKE03kkJGU/6Z51TVVcva6+di1cwygd7ul+8MIlX6enCxJosYhNiDLSwS/sbbyqbdYWW7N43
Vd1HF9zfmYZr0+AlgnWAypprxCJ/YDPKNcvy40bHslnYQH4XIkRjkPCpK+Y6W/KkpC6men/ncQTe
+SDfUuEsKf502Czaa29tdjE8gWnSPP+F/uHwbXMiGEpliVnLgo/RkUr/TCkhDSowV5H5ZU9rHFGa
x4qqFpGwxIly/buQe5QEAN6+F2/y4+1rZOMqK2wUrhN3fOq8UrVhvXJqaP/84v+DKhf+5FnqHZUS
JNGZBVzJ+Hmymm//FV7ZHWj8xJsX78UmR8IAOTdFegSPWNCD/4GFpSRZ9JPLHcyBKbTjR4PW+gQw
HuqYHzFajE8fg6XPY6kE1zMw2mHcZRHw4ao3Li6Umwqdh9w932fAigZ8Q6XEqeXjJEtyoyXD6tO5
JDL0q8d6RJPgAOJ8VjqnBtnodkw86y8bSTqmSDo7iaLbqFUgby4aVUI7VnuvSSf7kZy/JuwZbt76
JLl7yMpyIOz3jWGpB30oihTZ85CVZ/wgBGXI3md/ybw2Q7X2yrEV1V9WQPTRqUd/QmM/CMsdxLB+
50BVsZmoIdCWeigF/KPx2ONh3MDsvJzmYz1JmdV6s1kdvnxpwLttQKpy1f5ATGCfqvptqYawrtyu
yL5JaCu2Zjj506AVlwwHtpeuB6jJVXFESI12v8r3u3yXAveqwQWR05FW8Hgbkw8GbFPzSVWUZKHj
7M3eK5hMbT+lQSNQyse5jX79apWvplFNGuEH1G2jnqzmF0CB8vwNo2geBOfm20jzLfys4msRxzg2
KztIMAZ2jevR/ZwAY+eJtGzRGZ4E3f6rjlq48BFG59KnethYWBW9ar4qrEI3QfkpEQZMwrIaILN5
C/39qHV7bb3o255q9bHxD8gLYNGY5uRnOoEBK5CjGM9X8Jn+JQS6/Px6/S3Uo3jEQdNt65UAi4/N
BuMk57mMwqZxq6pvN/gia/Z/lmf3bUClkNlruC+BLJN3IncrdZ9/6ZjuS9AlsESLYYXwvhpMfqi0
MSbxsMwchiP+FP7RDSrJPHvX51ven43kD8oB5GWRX+Cs9Hqx/P4ZE9Cf1B970JmbpfsNxUpYQF5b
0/y07h5PLbs5cOkrMHvIQFp6SpOZVAfRULQLwNBEATAW4UWU1KrKCFFNBezfXlT2e7xCHNGP/gw2
pcIs9YB04mPFh7nRY0F5mdCsG/HNC7aU96Jx4EzJnFxOMhbBprbS4vco+BY0MF+0AOzfjsFa4bMv
F7ZFwtI7ftbBzWzSstakaVKHY5LFrg+ypbZYc6GyClsZ9Eb/WlyR0B7UlZ+FkOMQsTm5KYS36xw+
MGdoqRRiRbIZh4v0+JQmA1CPG8K2NHEIJp57MUNjnMMqGRZxBIHbn9pTHtiOQR6NxHQBIgmjyXNH
FKnaYnlm+MJOvwWFJCEl4JFAyesJKhD++D5DDMHVihPH3L7+My8B5FLrH8x44EK3O25srKhlGpVC
dcebWkIAWN857WZyUzB1rdvVbFJ6NcZzqYlUEG+asRmJl56Rn59qKGujMMkZADm4SftAs2maz5XC
+IoFYFPFqnFSxqb8Px3XIKTC7/wOp2EPLWzafYxHTqbQt1KXGHtmQXrtzQyYATMLVYnNQdUdSC2C
NCgBR2EF/vjZ0Cq0y6JaNmCgbMw3iBGmZgsXfV9qPCQQUD4Sj4MX0qmoHCTdyXan8OQXyj4szSWi
5U3XQEYfyCzrNJPOtHqWdranuRwpAygkPLhjItpoihjdA1XF4jw5SUgcTzskgz71f7Pg2IQz0Mfi
Tf3wMTt3hPAsHooK6JvS0Ei50CqL6KjJYZO5OY5ZxNO9wLVNv6Yi4KL4yOCR4DGgIhlhz6exAoAE
4PGsRyegocrUE9aZ5vFekYDsQNb/4fzUNFBraFM5zeytEWbE8bpG1HILFK3O0ast9vWPpkvHg/AH
6nXi5xwUtkVbJ4eyF7wPIpW8C1vlLmaFOBKJ+UG0i1i2qaORFt+IrBW6hzPHmQj3P17virNSxob/
UpBRWsLem8l+9Sv6XMBqZJZGOT8eIcAC3f1YGuesOtKT6Ob0ylx9LRwCKRD+lmL9O/m+uI2e0e9V
3oBYEl8rzeVjOWKn/8blMxNx/D5d9NxARfLDoQjuVpWfblFbfhElI0HbKPMvuNB/VDDhP0JwPBQD
6yCYP+p2Z2uXqv4G7FE/4hHK55AUdVRuvhW6wmNiixz5ZhCLz4wo55Bys/gXqbLL/j0Ft9VfN3O7
jL9hno+DvU5eqvhllt/rf3j14AxfonSV9xyu6hpZxlClJ0475prjV50c3lWQsNO+P/9aiU/jyqBq
1UdZGvkOuXfDN+gEtueztBNC2QZzPxaxB6/VdqptucB518/XxjaZvieDYeprrvax2/K69GFjmS+X
JWew4GP1rVuOAXK3u5g5MnfKWtFnRmKVLEZ+YxKTT7tvwXEpoYtxDXRPnyqlFHYwOMxOXmFn43f+
EtiorUNGRQskbNv0mUcHQwiOGVZwhrXRZeiUzsmxmKvJieiOJHgZpqbeuphE8TR+n64uui1+g1ya
H5DnqgY9A2WwuddF5nqTlgpP8uCRzA4cqLeaPZBBeeRLFP9hcYCjsv3DXH5268YFX48RmPTtlVOM
tpep1CrmhEV14pIQ5gdeSEfO7Cs3/8pdnaUC5fadOQhKQqUR7vnKgfAGkP8zenT6uf4wmNJ6pryY
l3mdTjIWO91auyj20G2Xf22EKKfhqljUY6CGO33fCn4yKe+NBOqBCCqa9az/Lbd14XMzX+/53uu/
63o/YiTqYA03sgMFkZ3BVC/aYcpsPI16RcDVe7Oe0dFoDrIlT2s8MlzfM4z3R7IKYaUnd4xpaZgE
FA0Pfp1bG+oh6kFOmIpLMTu9LZVFvHkNlH+fGN1qPTvKQqOlwJbx2zdO5Q6d413XuzlIT48fECDI
sb4NlMsgWrFRk0W7rHkKmKGXj9/9gQO5XtU2uUgXsBF/6TvHcW1LmMVDbNBfT8OJpbuT644aDH5q
rmANaH9AL8Uy2yVNdSoUzyqsGq9inv6tD6uqvbSjddCid9g7VpQm495G5ekqNvmtzaGXv746C5Fy
fFNWAC/gPtyP6gM1w18KoF7h8RM/aTIENITf/3iT8se/ZT7qCCONBGLxvtwHLgK49/l6BMq0eJml
FsYfOyx63Kkd+OdAVYvKtUrrbqgSePA2dX122etmbK9/Ii9Y1w5oNXs8/Gy1xhG74RDaekRhvc2/
w/IMymzXSvYEBwNUF+Boykjt6aKIaZfLpKgvxsD+ok1MXT8M5Kupb3UIUEdBZ5Si8fJz/J9h0MjZ
GtO3ATB4reH59TNkn+gwwnTuTICgyUtJ2dkF49JuUkBfzK0kcmSyq0eaNdWizhxi4Qkywu/xw0qg
P+9TyyYqIC/d9wiDm7q+2XixEMCsLXCvdAW6gC0NOr+4ej9NOILPbp7M/sAtHmPHK8dVJKaoKqBr
ZO0rpA859FcGRGubnEhI42O4zoFuqHTSwrSCYduvLVFs6H9QijIAG2QSFMtXaRlZxCva737b4la3
kJDCOTQl8cGp720z4ALKBjJVSg4swAMmVvnK/J0fnV0C83DoUiKdpmdfsVcw3t41AGsiJxJ0SVmV
sp2aZjC1wPBZ93lUUr3j2k4/US4hnglJofB4EcpCQN1oLkB7dq3trg0kIYuG9O4t7MTKHmf/J1MK
OhIeRhPqt+7Cy0Bl+jlnAwivgznrlyQ5JbzA+Ps7lD3IEW6jIqsacMp4o7TbUZOx+njHzRlDzbsq
Kf2A4QDqf1wNRpMxVhv+9MFgz8qE9+OHdoTksPQMaxlqELRG8qxsjZO3KLyfo5+7BHFMuRcOKr+w
buUwjwEhie5+in7etEjG0bjjBNwBKiUDxtCXdaQA5lXnHp8VGE62VARtxpD4i+pI6+2MJi2wKVFq
DUWGlDmAkYm68pzHikGdJ1IOCXM3i/STsywcthqmebiT7uARNYQmq9xoi2lXIk4ufPBjLdHVjitd
G5bMtZtgWviVmFbRkm7EmkTZ0aHt9EyasN5n0XXiBpFcR4K7I+m+XURz+Kz5Of8f2UVP1p6TdkCH
kD6UEy4cGge4cU99wnq9qyDRirubsrSzBzpb93YY5YgRY9I3vNL5TRX95RSlv4VVvBwA1pfNUZL7
3GES6LwSkyN4M6CsPvEi6R+UIUgv2cZShyx2qPzti0o4KyHr/iyk0dQa5d6rcMFk6DHOMeSmH+uO
gPFsO2hmsMUMUqzL8ZBOVYU/+9+Aw9tSB/80f/ip4vtfds156vcTC82fuom0fqUFdzdwpJFdCb6h
kFFo6Jcb7nqHypiDpBzLy/R3OFPXuUgoajNqdPf2+KkMJVovuTcd3SbY0CiqV79XsFQ41tZMwfIX
jTUVxEaKAvSkL5Ak87bSmKLfFlS4EJTh+TvxEeZ1rjgXNxrClrCTfrFj3W4824nwb4jv/Ni6wZm0
gac2m4iTNKF5QedDeVBXLL5Lj5eBnNtLxak4Q9HITRdHaneggypr95PWXpx6JKxKrPhIOPHMfosT
wyHBRs3gbxFSctMds1lN9RsXcptIG+ENeTtVH7UR/Hkj8GBH37n8TJAYJ/HiHvF+Nc7fsUN2UuZW
WrZsglBvYcgBXY612rFWk8RcqgWe0HTD0ElAQPJ2ytfGUmtAzw1mcmVznu2kQDp1JtniulAnvG9b
zT2MqRqOjoARtSVwQUD8GcZD0zdWLu+u4DVOHM4NJ0apDn1RRU4cXPknITUACeTW8u/zxHoaL72b
VRBL8bcUxvr8g1VCurKBOyqLhOf7GG/lZWFdIomECynauF1nA1waQF3HWXFpLTrk9mYDKznlewPf
yhaErs9goqDMtIwe+3AtczdN0zBty0ND5PjhQHwxr6xmrtO5cOFeq5tyFuFkG0Cjtan3d/Kucd75
TkwEnwGkXIGom06uWiwsfV0L7U+gzxbzYQUpRZNwrkFxJZRrKCnoD9cFbIeQ5qJS1Ly/vm87RCys
bgUSGr26WoQlHwp/sRk+1EUTXfeQUBUXyol+LE0dGqbtVTvUba44qi86Z5akuwhxXyWkPkrReqMo
3L6xN9Ow8VPhX5IT4BCMLeVvLf5Hnj+e0S/LCGZQiaC86m2NCX1P9MgHvYPDIqem5sE0SxAo6JzK
stPNnGELPfUdKX+vNU7qy8wbwAtN8M94xW02IpNNSSIXyzYUgBUxh244K7EalZJoeRoieRamXZSs
olkjHW2A9VId8sRl//Wb2f022IfyobG5/DD5Th+JeM1umSRHIJxZQW/+mTyElbp+3c+RRXB+Awew
LOXDYvmTQBNtmazm2Un78pb27gzOZPq3jT+AsUbsTOCFOu71hUFOg3RHUAY4Xv6NKesvUtcZxLFF
tJ77LjzZT4NfvRNmeMHq+BT4Xjt5WmCLRYnanvJS3pzkZCItujTWbuIRcKAJ+6I6W6rXhkNt/1tw
eth1/ldHqFtOgMGzCg8DyuBTHsDI9uPM2IbDJF5fdkiJcQy/AJOz/kZz/FhflYW9AafdEzsGaEMf
FqXk8oFTUK4Y3BsHWwS3dQchjfEFnOrGhRSKSv2mTmDnmSVFdaUKpWh8VnoHR1FN1/9IAFah3QnO
YfQbmfL2Xb0UcCaZGWpLaFn3aRENRnqIqbtRBaNB44Q5kvFz6Gie/aWlxZiYQFHuyQV0SEinmRMU
+TZn6xXnQ79ryAEMuRt014+L5Skmkqn52mceu7Q8BM0Wf6uOi64RHg/lcwuxeUv/Ok8JArMJgjQE
62EP5IZfSpXsoIaKDH/Db//w75Y7f9UAdl4/ECRwVoaqDhk8s0C5VemHdZuTq3KfBV4umypKp/SH
FlwUakstjbq9d/893CwXr/D5QnBuf52K6SGd6fYEsSoivCtJlB0gteNFLvYL12Nsw+aMpCDPRq4c
XDFfYDzokq/JHFL/EWyeoO9sZ2wffF+2G6RHHdP4VqhUO9HTWi7vkC8AayuR5xs5HAVtp7N/88DY
wjPUtgYAql3bjVe/ZyizU+N8LCPowrjFaHYtwmPzFyWYuNFTfWEaqcs6cuafabtP49qjd4QP/0+/
9zqpcuG/9RfJDhpiGjsG/XYVj6/cIVpy+d6fCt4DF/Kn0oaZZSf1F/4cXWhgjo3+Gm7cK3NokiMO
dJET12zFm1aDoocbYAp9MqmmAfOEfnYywYo4H0OyRUYNvKBy7Y14QCyDrA943UZhwLuyXu9HHS8G
RmbnzoJUohApcNsfBKnJwLT9z8y8hQb6+mGjXAhvxTeyFfq/3SSJEnQXV09LFnFbwOjtUSXJRzQ/
Czj3rh/rSjQC2xDi1r++RO5Pip94L2FtSyjg9yz/ZIepH5Zczb5RpJDg0wa4p0R0R5j0bojJvrya
PGHC7/WqpkzL5rSOMM3v9EvLtoQDKe2z9OjkjDBdsrs5+69HR++R7OnjQgwzT2P2beNmRnK+Ybc3
QzYFeAq6YTqLQcM9fp88/KjNVmGYixuMGYJNqcQct5pRuJEjX0YgLxMIKxI8hLP2K0+NRdse8d1M
DmF4K09mcFMPv/GOSYzK5GUnXDEO1XKgCk50NtkjwvApAmyjDZsYaT9/dfF7VIWmD0sRIKL/xZpa
t0bX5hOS2My0j8luvc4ARsOIqoJmLtJmyIWyEDs3vZhef/k4QHdOiQinGHE3f8o7Gl2fe5ulQp7c
MxMw1KiyOgxphijByg+YUDyvTq9ZrvX7dA+LA7YTa3B3g+Fq2+x+sqSxr9tM2Y8YJoXPXgMiireQ
gJQSdZx8IQgQcYIk0p5zYrXUZk8vLhTgkCQa95wsFnNcitGhiBCCevDeHVl06gLeXr7OiJSjrIh6
bn6H0yDX7jKNklWNcW6nzcGwgIVIQXRnuJrzzsyINQeeEF3IDKgZ45tOnTvHWtWuhuZXhaVZGHmD
4ouObg/BYAPqQsY0GEHo/8dXTh56MCA4t3MWizVT+NPTsYslYgGRDiz1KaYXF6fldPZRX+QxDUlF
PjiQUtfzl5VIfAS6jmNZDgJsrl39iWaw1vSQKCdskZglvNfqAX47PkwuvcM48auZKK9tqOzzdcl1
p9IW+U9HQfv5Dluq1wuKobxA9NynEl684ELtPREite72ajTnozKYSK5YxnRPToeciFWkT0Rxp1o3
02153RXHleFf3mI+ZQsZSdqom7zD2M6h21dkFDq8YDISG5yYF/aRnzEu2k5CJYrtM/KpZ59b7bOF
+HbzgvyKqojjioxkk+mjB7YDAxYt0fIsPH1ePr/fgDQCuAKzcM7My53hGtjY6eEQ/zTd9ik92+lT
m8I8/WWKQVgPqqprgxbKlKJx59VWUquqdd8U21D1PdqDReLsCCOCA2CTz/XVI7jrzjzDJNRr1Hnf
csaub4cHXILhjoUpim9JJ6ojTFfsHk2I4fRUxXHeYySdYSStyVNw/DAkPDU8QVr5ZIS8klHAnELC
Ofl8Ewik4GpmVBdjbiCc9EyerA+kmzIO5ZpPU4Sh/OJxE87/aelLWAhZutWqnCP8OcAsl8prhh0v
+/qtOuy72XBl8ZtkIObtQEXFq5MSOxsNwFb+RoIOP9Fm51hY6YKGpL3FWm6hcz3QMIlEkkzv3BCR
SeOgj/sWvtZ8EHyh+ZtS91FWyr5mYGdM+SbVFTxlcQnbmtjrVGE1OlVbttQG+Cet7Be8f+3t1m84
vNbE59ZuA60rXAPe5/x8LEEhFkjABBhBp9zIgLtNrhmh2GXJF/NFU0B2xHjD1x02HE12hq2QXeJ9
S1uVMhy74iDmwJndIjt0kSmrPtO9F4gkFVla3VfsHti4ATt9t2OjH9lOmSbO1PrRB+0gLszpUZPr
FscclgKrebmSPB7uDbc0xa9gGdPbnz64V56q4oh/7c0YXlVLbkbfJkF3OGUWarhumxdiL7xfTS11
Zcdo/Vg+FyVc+kuLHJgqcSHbQbLYi35CHEZeG475ouyWJKjTjmc0imnQ5rSXeRsAXcmUSw9gbHDh
tPoS6+aUO1b+B/hhOpTfQkf/bYk5PwBucU8bzQMwsbpziMLLuPJp9gH8fbXmUBK5eB2W45i+qmyb
1oo459E1BXw9jo6e7BMw3mGHogl7DC9Bn33t5BB4RqkVVs1GCwu78a0HH9KvS19cjNVH+hxSubwv
9fLo7qbQHGS/73G92GSc3rwre3j8p0tTRBiYI7dLCgrnO2YYc9COO6xycjuF3pjs0ri6JnYS8jsc
2Bqe2+0aHZXmPvYdpJGERgFy3a/AhZ/NuV1oikU5UPxCJ6bYHDxTjxSvEQWehw/xzsvEeLJVh+hj
c5gtf9rj/cvhWRaiIWBbQjL1fj6CSsqJ5p+r+hhWjkxj4ydTpjG2gR73ByB5KogonttXBYClxb7D
RCbf/97iJVXDDRCNxDtG9vp5c+LEXryAg6Ed1cs+s8XsuzxAhGJKq6TpCtEtBLU7/jpqnxjpgRL2
axp2DY/xN/ztZxTOdHc6unmupW2FIyu2wsVZxFkbBJzDZf87s3rYzhluviTQqsQLnWHHmR25Ygrx
osRvIKKPdRUDavWRmFR5UqUT8VsQ7V9ijwZ3FuoxmoyC2bOYhG5NlNWXH2/Y8WP8F40ih2Iq028L
W5IczfR1ap0hpFK8VuKuB8HspOPzsjnwVEKFrj2AunvMvVNsiQQigdGsD68bWeP4mOf7aYdPlNpX
3w/tXM2R0y3h3wMqYaNBbcqktsafeA1YtqkYUtN4i9GTS7VXBEFW4TN+NVn0hv5OGPnOURWviKhV
JGkxKQCf1xISWTqp6niA5rZBAqs+aol7aPFw1eHyd4Sx2+NnVvcQDhseqMeYtyDuuL2p4wKU+Z2P
DO022mChujGE6NR00IMBKyCdIIVGxCsYLXTH3CcSw2ZihcS9HK+Xeq6CC7fJK8xOTnZLuSOyR00o
ZX2IAS4bg0LHG8Lh9Vj6gjW2k+dXj16+Xy9+jBN6HTon0S8jV6GhgFfRWE5BUuHBXiK7d8K+mtjq
+1ZYZtXMgWh9qDnquloi8BRDcqrLjaK2Hmci/EWJTNqzLEl6m6Kj8IICkE0Iqg1A+rUDeA2pbgU2
PIPYEujdpOq8pqrZ48ra0Jwkh9GhICqqfsv9a8euXL58fnsagc6lCRsB8qX8rM/q/E3H4zKAhdSK
AdHmyVIYCHvuRCtPH4uZDmDNaAzrwy36dGSwQraeknk1vevnL+cEtA9yI1CYT6Xu9o+m5wZ9oMm3
Dna03uqf5LsV/xwCVS8laWbGMiW48+CZNf69fsNY1MzXYR71+ph86zu+6Hb0GKRae+RcR3UK4lhF
bqqfT3HUtKV+J2cb/kIjCgerL9e3om/rPaR+fxf2SHRxXzis3wD/BV1ifFcvy7YcM2yzVZ2sprj8
b8YNv0r4fd16E+1+CrSMtrtPMLw2opwP3lWfXOXiRoW/ON/5PQ64PX7CV9ueeBwnbwSCkvdMFLOT
KquhCov6Z+JEiTs6bYyfOFCu4XTZ/c1qRg2mnUFZa3mmQ1wEVzqTqrmKiqKOqA6zn1wzdYLDTjKU
TP3X9U4tip3+f6IsNiE6BKTQiThAQM0uG300HSOZwNhjPdaPcfdBH3++LiWd+o/YrNlj47VVDfi/
rxnIEQRaAeM/cjmY27neO0ZduJAgWVyv+dDqLUWyw1XR99geaqTrxj4ejAHHrrtn6QnyaPcXl9dJ
vObHdPtmjd507wB1DyWsxUMQonEDt9nMhZUUbPfhDSiWZnBHNr20xnb8pxWvfOr3RGf4rk2+IHYA
kdP7tYlicUJa6u+qi088+RaduO5TyXgFaFMmMmVJgDInl7bPCdhV+2mJg+Mrc81FIPuWlf0ONPPC
5LSPGS1zifuMo6yyTzMZXJTzEW6vVc36PlnpHlxdNoJ7aWnyIvto3GTrGkgd3MFHu4Q85eLZ6XLB
WU8vkfUN07+Cw1Q8+/vQUXLzynvu4J1vjylvRx1t6gVZWUQ8MMu4m5Hzz9PXm+fDo4h/b5ok4tGK
gN1o2ESf20U2JP/amKxDIFNrsi8C/yLRzCeksfb90rSWnYLKZviM2m9oFx/eMy54o+Jgs9wiQp7d
i2BU4qXcfcs/Xkhf2d6TS9x/khbLEVuDDnP6x7fy1jS43DutOXuIlOhveJ7kEBZCa9lph7O2YeVg
TKGpq2bGRSLNwTnZvCH0tZesSEatcvg+YKoRtGeOLI12j6sjW8+4sZ+kSbmkdvk3VhT3cqLDe70q
4iRMzmGCbq0iXHu8NMlCztaHpCXIWSJqLe28AQM88qFPFMxiSlrZ5bdalI9SJHXmhNUnYNG+FUwp
e2qExz0Gw8sS/3pLPAOpNgWwrLC6VfhjrVkGfj0sp0WTGXyz1QeyO4cLvmjoC0NdH64ledqo/FeJ
PY6i1hVMs4cTqNuHNy8fCUTmWU7jgveGv55AtBHc79UGj3iTvfELl6wDrJfwT3y1haV/uoVBd245
rdRUy3EJ25UvGATAvpBZpAPU2j5Al3aC7+/p+UwbJJMuPzWFaE4GIpffZVCEtM86XEm9/qzpmkZA
QSIO7dTCt5/baTvCSJJtEnzNNmQ28spzpiYkmAgZK/YiFAPyKHBb8hDcJydYVYRvVDGZxSeaTmtw
sHHmVsA3W04R8W1SmNeyXJFwu5+SnEZw7d6iFKtzcxZ4g6xqeZLgTlhZk2UH30zpXwFxTv66pb69
3FLmz8dNjYNm+mUh8KzrGblszaOR3zlhTO/FARPeY9/Sv3LCLUXrpBnTpHL+0/Nsf4b9EAVixL1W
rbvVeHXTNLxQMC7+NNLHPMgQmHrHAQsjJNzFqwcYdLR5fXSsFF/zwBS8IyRcZsFZwQnEing7vbwj
xUlDLLQjssYl4unJVoWkClydC++I0tljoNlMsJipWG/ZlVEsaKti19dAgsCMc48i9lNKSsNxDGI0
SbT9hPFC0VGolptR1jwjyv+JrdeBURDoj+pNYuRVSv9FVR/pyj/fr76tsrxB4qbZPAPssG1gfQSt
NbYlLNhuwjQj5KHDj8Ens6wkZRfsZ3JT1DVg25LX1wHKtNPY9GtSrMk026KnE3GlxLI6wnPj+Uus
JacePVaJbrg9yAbUB5uWtG0IpQ2eN3z154KtuBY5e5bfvZxZUMg8CbUKP5stq/EetSXyKie254/o
fXHRO6O2dJjkT1b3SpCOuSArvuO9trZXfrkmEBSTnY6X4mhb1+ejuTEoAN2vCCeIaoiElEdhmtg6
56/sheFpi+FvdtzzCyk8r8g3BeYG12VSNaQ3Osfjfj1B/JnnFYz7d9xSuNFkq8hoIoheDfJlq1UP
iz6pt2n1lPrOaz/+iO9OCx0SWNdHO2YfuhQavLDJS+pv2LgmmE3aBT1nVj/6B6eMDZ7URcuEItOu
1jNlH0knc1TQvLtW9SIO6CVKW1ZrFswKzP5O6JxUfUTjnIqzFNA/qgA7G5Zzk9yazq+f8NCDUDUI
XMjPlnhe7Fti6W6fUl2YRQytftIjR97+5cogmtF45ZCDRXqHmdpjvsq1f4r6G1LC8tZzA32aj3XD
Cep1ZEXikJF/1fXVVF6cY+/JKPokYPtCrDEBznO840ORIzAih0lPaGPRaG63ya4A7Jt+GLWf2g+9
eFiSIyDJggvco8tR0b+6YGSuFVzepFiqpKM/Cf+GVKpb3AzVlbQaMQzwT7tnwTGaEsvIznbFDFgs
X62TzvO2uWN00e/AzqpFzzAAt1VXblRjAw3UnZ+gX1qvb80lFZSjf/grAoBp85nmpJ+vJ70nnivq
BqUzQHX0qhg7MnVcl5/Xkab6zDj6o3Jr84Xmza7bx+wam320oDbgqqtT6gffm1uwiYKCQ34U7ztt
nzpzDPZWbP8R7MDy0a129EL6rzwQjCnWP33miewlUfGCzOzJH+MQsZtyQnHH4w6BgZTf7c0+eDof
evEU4DQmuV3pLdNWmERdkb2f01BvFzNvlTrwwLurpLYYib86TsEIPeeD2k2Qaq2iqHGU9WnsMTsR
FgrH4bljuGYW7tJJHCp4bY5JRZS8KX6utDO3W1amMpFJgNqyoz0mNc3MEfwfr/JRV4eAPkO4u/Fs
eE9xhkkziOcgxzhu1K52evsJan2WZEtL02K6HYrGSJkWsuRMD3gF5BLWqfNGYz6JJc1rgcu+1x4L
9Pkugems4o/8uHofPea88pbXg28nT8/93T7dejBhrAKCvonA3GPwdN34iPJLux7mwFm9jAbCKjnL
07GDcx651ZzWJbytOKgXgWXqJ/HmoCIPb8zFVMGF8X/ydp1Xc9tWsqdns48ZQ0/QywKKxNfhScXK
rNmnOICRfnQD4j9bLGNw6ki9yS2/BNX2Ady1O72y61S1snLH4BHQw4tUjShT/FaeqxJedRKmd4gQ
EwfuPEQBKkUhHuDe+QEYdlVhqL7jp5Ra3LjfdLLe4mnPHR26Jn5OkJ00PDsw6t1Rk/1ZxpfmpXY4
AxOHDizxMMOu78agEQy/oij2G3h0aer7iOAN2VZVGF7rbjpsrqRXAW5GohU/c1DVCNzdtI8KF8UF
iPE2IzbLINiTLv5ONtRMu1NZKizjmzCSRQYxmkcsdTCxiNJQOfb/MjA7EEnp2rAWHeSsFF3+Ew/K
d2vDg77d5LF50RtwhpZByFytIIepzAct5J2l1P4u/aE29iX6svlDoyRXayh/QSWtgIeU2dN9MD7Z
Tw1oQLE8W+hVfhubzHu8VQZMIiMjmTEUOYCeSC7Y+j+BeND0oDATurR32egBLc0oRJdN4lQ7Iyea
n7dfPKZ2ntdn8fxOY9Rqtjtc2UnbvGI5txKakCpXC8Qa60MDPaihDJaED2OG52o1UtGsi0Ka65xu
YRAor0BGKyrEB8zunE5IBueO3hbo6a7CxwjYsvCt96W/m61gVOytlFU+yUbnS9v3mTsOgBh0badM
uzgqhHYPSUukLQVtSIgv/gJYRtwDyd5KhCjH7HneyFuU9Doc/JMjdUeXDz6P1VFXajIpc9kqjOGl
fxKvdiMi4jyli49wH9HcdIOikY2kjBSfNlF1hFuRtROmt1eDqe7Nxvh7W3WecRBfNrnB1LTJUYZB
lD00k6YIt3nw0DLHftjLg7CfCkjG8vuoR6QhCBS+4zChsaLU/t6F/41KsZQnLsxqXydDRZSPciZW
SrkFRXdQSgoZ0MNFWhEENtF/JiNhbZNhLbmO1wdH0qvL5QbVga+CC8rd1VINblsi7ePxjQMUxlFC
UFkwhJLdPVsDos5p8i6MRCAuM3Zgn+uhCd2eGcfGlxZMLE9E+1C2CdcKw/aLy0kHl7MV5w5/7UOM
YYsIKGBzKw5J7BTKy6tASRtuszK3ESm0tqVcdbEW/75S1g0bFnM8BdVnK6UHKUIBZHOzzHVTawoJ
KQX2pgK38y+QiOmVxlbMNXEftfk5AnxJAikl5OL/1DBIP+sEanp3a7HmVROIZgfiV6szNYYze/HW
3YG9mEU5LV6AewhsIWLmyFQMNpo/RnhHMKmHKKfWSv31aKwUEj71J/iAS1tyM/ylz5vd0nQ8iL8N
q+Z2gtpvgYpCzvK2FPQMv3E17BBBMRfVI2cqBKPgXUZzh5UsVtKu1uKd/wIhYs9SkeBReDyw/cFW
tJ6fC7LnodU9TFXKUBTEsY6ub10oHsG9cq1dKx2rSQV5QENNOuEakL9yySasLnjsMAnCf4GuDBix
IFy21mnMvOO2vbAX0d+AdZBEvNQTGVGLAIeTnGsiPkhSx+ImaXqOGWFRge5dURQC0PXs+XBiJicr
sM+iXenfhKacD2z/77j/hwKIwZ0C660BVuMrbKwRSBqt4pBYFxbwSrfTmcu+pw/00auuf1r7c9s8
utcLA3J9NEDFBcT8hA49QAQryB5ER6XzYoKQ85JdIuQlbXZ2svVSorEY/VQzXbWbzKeIUeOqocoZ
csivtodN27BiA8uJ9x+CsZlwVMtbele4HGTjMrSNzTI6nQlSgiQiSV81CZ/rdf/QBv84OpEij9Ah
/NniLqttOLdJateLJ2vgPDhaKQmu7XpwPr5YH8QOwXqD3ocXGxHhbQF8kZSCCo7ePKnLNmlT7oCA
/NUAHrGYie6sRT8qyk3E51mjrhx1e7P8A0miXfmGq5WZTS0QdUIYPG5STKSCugoInAanBxIjbQuz
1K2gRetWNagMhf5rR5ZUzI5xfYwrTraWCb9jDzKkxU1sew1i/XzRpbaDyyPrI09lpr0htC5f/HiJ
FOs3kKERZZbCSUQ3y1+2l7gTjLS9kFpD/iB1+Bqgc4iRoYK28bEEcPvsSTYuVGbB1B/lJ07jYJAo
byHgNjyf1ot4QP4LU4WqNfgrA7IPslBd/kciNbZo1ihDpoAXN3AO/eC4htsTGrtyNfCEUeKWQs7f
KXaNaVV6jaDbB9QqEIYLOTaeCLZrLuhsz1tMnMkbhO50EDh22XzY+Q9l2knuG/ZK+MWr2MjGOzqa
nVmKG7uIegsTpvSW9MP2VYLjT8+K5d/1nY6VpF7316qid9pTefM1iC7XncUGHaBjjKFpXpj1tRx2
0LiNXCrgkSvkBbmq926wQdcGuY5GPl9dGj1aPIM6N6GaTK8UJ1Knqknw9tCQwApw3DdFPhYm9nj5
Ufq4/fZ/L9TWwcosMhsn+zJvHCKVOCRufNAeTUAVqRDpsrIi7u6riTnbBr96h3AyV7p1oWHqpoAo
KrqqOzOS3+jOxPwLrJh+jHT9FfzeIm1ihX3sKOLwXbc+Y3bh+TdYAU+fgM2+gHAG9JlojW06LH/R
NXX/0YHXhQrGHknLDSNjPMXpLPKHIHz3TpRHzeuIETT3tff/xfGN4NmZXMjWYXKypXUlZVENNeob
iGYB2pJMHacluIf+ud6QxEknZPYtSshhakjNbhKoQxIovOH8AnzHz2JWB2j4CDPgU0IYP237VsvH
TipFU0Sfj6VKSPEHFIfK9HvfrEJFOh2kWQ2u29sTyf1q/W7uJKNIVjTYsSY3Z/Ocz7fMfTINnPzj
HlOojlLRXQm7PDYKdgv2lnXK9dAuegKJ3kRQo+qsF7Wh0e4S4tcFR9ENpWMFFewGMW+C5Hq5MUHu
toMvSucPeiVj9wLYEGnozBe4bzJdOelkOSwfWQOuZrL4B2+ZPpmveQpVyJimc6WBTXyxughzzw7I
z7MjC6klApEM6vZjKpaZdRegEjLc7wgy9l8PZWuWdfc0VCgZj4QoqUCIXEHkcLudfc+Cgrnb8N23
Mu2Osszi+/+/fSxR02U4sfFeRBEo46dxhx3ldZJmgdfl8G6G5Q8cjwV+EfJrYHGBeNDt3i++hEkZ
CvN1d/q4zXfjW9jKeHrjRYUWvHaeeHblReyBRpMpT3R19D79HXNXfD/tB+kUPbKSDxUlbfqy3Ppq
pqz6QvFNGcmz/upAuXMjT6irA96CIFXJBMMfW4X6C3SMpWo/P+yFMc2FNqNltkX3pxI9KUQQTUnk
iT+SoEE8TR1C+h2bDrvFARDpu2oJMGiOrLsALwSvJFtoMvRZnkuMYXYWlDrvkYEQr5/QOWhNNlax
51cMVO1WiEtzH4pXanlQ4xUpohX1EcpBkV/7HOi6glbbRSPHHuZKWbROnNjlefyLjJadaojfdtjc
xmXbCXkFx6Uqt0go6cV3Dn2Xd+fgW+YRLGYTPD8A8aJYSEjOCB/HnnDJ+Xeb/Rltjn6QxJOjXsD0
NHFScQpyfSkA8s02YlCIxMOaSQOOulJSEFvTUx8nlscuJ+jAucdkoom2ybx4NjNOPlMPIvD0i2e1
OT8ywHGfXKE7jtm+Qi3e8ltWoYoI8gNzLFVxvmS3r1gIIH8/eaayqrn3UbdMWXku1dj0zdALjh/1
FWJA8KHg2aYXWwzTgdt4zxnAxD/W/exp9t8l0mhATK4IBHCvdV5sKWFl8dojtgFMi9gBCAD3OeOb
QJFqViTBRE86sivOrOnB3OSMNoyf6zjEyS6RzTyeYSLLNKas9GJu6LL8nQmQeK0SSeOJX7u9tcSz
6Rb0cPqhQZCPqpAfEJriNtm+g3T8pHHzXIv5kbOeULIvfhmWX69k9UwhFRYvWKkkY8QB8+8rDh2q
mNM1ZPwoyIMRJEMLmsMk5VUKNiwqZAUiY4xv6CxtuF+9JwT0AaMQ9l3RM3j41oR0K44dCveTB3+h
JupKztKGk+zMviMZ56mAlu80/h9FWyhQ3nk2eGy6uiL1rNgFCGAcIeejXDU0TLrvegXi7Nw0/27P
UF84ZgumzgKEwZzx2iJ1yAcQ78ba/V74L7hJdBQnvgCTu7gNqfeJkKfldkBSHsH4ovwNPROPP79Z
heVcWliMcFfe0QeRzmkjLrMx7db+Wogn03txk1yaHEhwn1YAbWjutT/xHL8lEgtJFcF0WctlYA8+
9uJOo4BUAm8XlrqQnf72S9TnmCWmBSM9VihUQVBbl1oJGErHM12m+ASV3zVaBPwhwX4XUUH6kdIo
2vJx/pXSZseSt29eMaQgStranVDq4SyhIPpR+n64Y80zJa6doaW8oOpWKdksSB6XEu7S7/CmAvtB
AJptsUp0oTIuoco6qY3lxYYG+VpG60kxg1BrCv44e56tCMF80sx6RaZIQ2HxsdvOBa/SqPFHwcAf
0lbz+BXYkwdTmXgtjUuYKH/l0xYdYR+zwMY+QXJhtDUxClXSGw3BQXTSRixnyx5yB3/2OE1BN3/A
Alg3Vnrj2xRthAoX2uR3znYOiHY/dvNnrY/X3OOb8LuWLCjx/xyDYFSpTyMKf5hIxNWpED+/FDPJ
ZoiStEbq0gU0zHjYrrKew9N9xgC3Y4PQu3w4S19sWBFx+UXpef/6tu3YwQ1L57w0FBS5/Kfb34+f
sM+Kvy+B+AtVA9CmTxcjYDOrEdkB71QilX+/y/XdzbtPjtKZbbry7+kJo2wgJYph9ntpuy9rSaKn
kf75uDSOVJUmvn2BVkHgGnizebg4MIpMrKeZs6w4rc9kCtJFuZFmbnvotcOU+hZnj9pv7DyAeydz
9cCxxoWiHmFatxSfRtRMlwYB5ndH1U9Xf2IKdH83tLezk7a5gVSEiotutjmUUVnLEbEAWhXfsLQb
GD7vVhM79Gm10/UP9Va0gjI9aAOg+A1EdMCntjSNl1gH87+qQbHFZ/bEQAPIznTXmdLwQ4E9eSyg
bDtwtCsTxXj+dAjQgvrLv6A96kJHBP5FD4nzxSZn0gr8zU1umC/nYqPoVzq2aMK1IzNi5o72qPPd
kjbRwlhF2kfrNH14sSHvlhffccZm8il9cSqKbA0cC0Qi/4gGiDJiHITEqvr9/U/2/6MzJGCMc41n
3Ggpl4A1WSbp0pIFNYzNjfG3+8kpgQN0YqgO4xEuKoqsnNTw4K9LArmX5aIsXxj5kowByGH0JQHR
IyjwMiOGVK/A6U838xBfkyLyO8kHsvVIScAoGLu3foYOc2chgzxhA5EXI449YNk3S/5tyQYYv/r3
B6Hu97xC7BY/wYQrKJKVeGITWAZCB74BNqpX8mxzKK9Z+iItERQFX+8njA+atsOHpj2XmJ2WK3W0
Sa8yD3Xlqe8oMRHAml5cAOaCF3oQSq7CQzQemB8IKcwI0rNgGXOTXB2+hyKFZwgyfDi7HjT7hBdi
NT9gP+/YI6jecZA3EcGccRrMujNdWVkkQwrfaxNr9kE3EdAR22LNa75lIWWjr/MZWJz9q8djQSu8
bShNWiY1qNJD3k5Get5W8HByBFGal2EOmOo2WncUcAUZKrfUSPoSKo9XLtgmgVAyiHcAh1TiA939
TAdffPiFIGWuoL9ngYNdeZVJB9nUM+BdwjSFdsbn+VAG8ZTmJw0GI1Kyzt+fz/nhgjOEm+GuylBS
PynwEBb/rBc/0ZX2IHO6n7P8mSCoYlUi2PMokaEx5RqUQrZs1PHVGVPFnir5tkLRauzI5SwcMjWi
vezWlqeVVtVgPbFcERp3pEtvS/I0YtJvqIcJFRs2nh2YEoGd0S8VqXvBWDU48WqpVHHtov9Tnj7z
s/AmKAb5UNxhJeD25b9prMXfIPZN4gPrZ0qZ4glfRxPE8z6Jxa76KUep4bIC/o2vu5MQoIe4nj6G
7E7y9rcxH2Af6apCQLVmwW6edF/IYP9pc7UGbo6d9DRbRBjbVcT2fpUBe0EmPubBFvyt1I0wFWv/
7UL8zxqX0OB3xl28G/QkHxx2zWOIw+jE+rqlH9URJ+Xy+nZiodCMQIpTnjYILOYoiN8h8VjbHN6F
49TgSEVmpmmZ5lfSa38Dv1iQCyYQL+yd/MQPmgG3cJPwTUGxPBcK/GM+YCjhV124wi3d19QDZqDU
jyVcrAqmUwIKICs/1jMb0t2W8/uWQhM4LdnmPoE51Xuy12wPORXrB0wEWMOkEOR+C65QAs3z38Lb
qKjAVGqG3GCrAd/5CdNNtIQ6aPj2lReoTeY/5DIQhCPqLTes0bW2Iwgl1bTBY+sPK6X1sRy6ZlE5
/hAVthw/h+k5aoDYHmlRTzcVayiqugUI2X4DMKF7eLJFwS43XxC88NyBbhuPMkGlsAA063s7QNZw
ZWlv81XGiVgmX0YUkeCaG/NqSRY2/sEgLBTEAKwOlqsn0+IRjomCRkOM/YITGgc9ldtWCMa0gfcG
tUad1zizacbPbWDgrJh/9FlK1k/6ZuI/owXOB7K9by6P9YeBNGNg3j7YjKdc4k2A0D7PmvltvcYU
MbrasaULVn3DsVfv0QRgoY7+nOmPDWbXKhUYg+V40lA5Ro/vkuT7YN2LVzCTfBBFPO3OjZctvaw8
+cG4ioGdEHjw8NSSBo/Jh7SGitfWg/+JGOmQYSxVcEzHLybjKpj6r/4ja4hW/t5BPlZGq+Qtk0K1
3aXRcwRSyhruxvx8ixXEbjDxe1p1qBk2Ra1RB8BEUgJNf+InWHFwRnVi0Hr1T5Lot6WGDFKdL59f
7mcq3sMibW93uVXlUDXIpOjZxfgBGIDOYTTZORF2gtCytXNBrP9XJqfz3lPWZNRD2tj3XWRkcuGp
tEtzAYMKUn6iw470jJBcpBdC0brZetfgvBWJqTo17Q/ZCz9R+NjId1U9kFdhWElkkkxfVJU+jSHk
sdhqLxdPW4XnicAgpQcOsAxCxDi7HF5aWIdTr9/PV2SeuG3MUA1Uh2eZpEwtvWBgZiS+v/cViV7Z
Ob1C7HSSqij/i+KFxaRrwGhXZSVkvBTqqynI2PP3/MmhoWIa35EuWkCWDGo5A4EQTyd0kSKVACp8
h2RivUCyi3wXqwlCs//iW0iH7jeh8MJcgn8av/g6xzI/6UXElniywPe2qQZ82jtAl6yc4TGCS0E6
v9Jgfpp9/q9j+6XK6LDjT7A3K0KT808ecgmomcjCyYKslgTCB6Z9L97YG1ZIIEhysnQ7k5MMAjKa
3LxIXqE+ugcoaxGQcs6Xqa2ZFtcCxSD4UvSHd0mAMg7aiByUqZ/gMqazP921ZaGsgvlfwX0bET+6
bn/FUbNOlu5jCepfKqToQFnBuRrbN7XD9ePsF7jJQZ7jiqyvwjJ5T9ohDVx1uXb8FZrDr0oWAumw
xd0yKIuILaqYnfOKh4lWBxky/TKUQsyvcQG7D7qxuaT57kX0bwIh94q6MDJK0TkuOmfRbgnxfayh
0TCKIBLKkg/Cg6+zywDkU1r3cMFcUwN3A9EVqUg6n6l418gTIEStS21mfn5i+/rxql5WjZ3kk0N2
UcTQkphs0WJ1kAZ5f5Ze1p7vFA4OuV5cP6LU1TX0vggWF7BLvN9mNcWcxtiOn0K9lmWp0EYTonYU
uGMFnvLtePgNMhA804wntykQja89wSPyj4xD9XEZeyHJPnCQOfpvDmGnLkI8AJCifIjZicJr9mQG
VOfaM7OlWS+TMwrWamaKW1rGCuw766dJdxiasCaaYd90X9TqG3wt8iavBYJZjMji7fsQB5QZsKOI
El95BY29ZWwA7KzZ9kP1tjZce2CEu/qfsk6Si/DJYLxdOW2QCPKJ0aI1EMwBrecVUBhPYW68DA3Z
wcAoP1Qx+tOeLRUmH4VrR1Dtoqjt0ANQaaBMDMXduEDeBzNLsg+yqOrBlHUea6bOe5z5unWzdUU3
SDbc3cDJSA1Zu+CkhP0seWUKdF2Sot6QVIpTF2EVwESY5NgKmLGAMSTunSKUk9vQPyloNC6vCnif
G3pHklBoPtYBppWMrgnftZPKLD1pU/mlV4e7RcgGUfmyfY+poK/ZoYXeSjuIZ5XwuuWjJKHp6GqL
4rrsMxMfcN0IBWEx1kABEXipkTRPF4KKT94r2qsyIMBrToB+2PcDgDEIT5e7h5bOyiXTpY59YxNd
/qJZtKa5EqVIDJd2ximWLF+L0pOJehvZWSpjY+X7GcQMbK/yKFmCmd7Q55cu+/41qq4YOxk1pC1G
VYDSlvvsx8rWr9/WCeU4kx2En8CHlpyzc791b0wEkvsFUxqsdVm+QKRQSyZBV76spf/2M9jwMpQF
Xxl/CBqBCyM45X2fJWnhZAm46hOf/8Rvx+Meo8Aztf0nTFEJgChiXvZmFzgmu97cDDjKfDZLHIBS
YyC4Jzv36Rmp0mlwLA1hBmNnvU+53W/4J3zdq5Um676ZaCioJNYF5Xq7xRZfpqcRTuBVkaIWAkGG
i2y7/AmXwPuZ5bVkcWyXZXeynnwYjbSQIBxoQOKEy8v2p95Yc76HCTq1ujD1XhlUXV+smR4jSbhx
wOFZKyk/fB0+AK/fCqRroh/A5KODErDL+2T0s5VLoJ3AY6kMUDYUopoeF5xe8m+yQI+cccnpY3zZ
m+dzVDBe1kCv+1mJlnK3PllDAoBhq7TBINK3L8kP1WLT97ivY77xysWOmjR22XSFEDwzYeFPXde6
CDoKqbML/l3E+pI+2t6K+xD+R6308PU4c3MQA7vwhvl9raU+KaoyyHOWTYXVExypMFli9ojl0lzy
dgI8Lt8NY6fQ4Ok0TtcHss5IAdM5EJdQBrei/T9JhGJTD/DtQN0nocdd1tkr+ot59AegcfteLlGy
+x7840mh45BdHidt/zyx2G8OBvwBPub0TcD4fGo38P2D2oo3fwhNzSuJ96/AUf2hWU8S/EAx5OXY
D3lUcHcG9xzWo36Xi6E7alz/sKf1yMHeJz+/KOIk5uiCjOo9eJAgPbQ9TU6Id9Pwu1xLAWa6omF/
vPwFBIk0AC+WGEXtaVlhwc7viv34qAabCItNInI4t9iw/Rpxwa9SltskkQK9x6W/SSv+4Oq9CFoQ
HaTZH14PQQJgtgj3uK0ev3edVXANDHcHtbkqiIdoS6ANMH3KKS4Xrfrh8lFw3RYL7f8kikKmGm3i
cO4/zDWiebgWMEdX/ajb+NTPo0AbDkcf69GBdeJGKQl2M9Tfz42nD1K1SWqiDfxL1jAqM5BGQdvV
sdknpetxXXdhVmoR5J75U6cjLwg0C4IEuiOGI4XHMc+akzzx/DCwZHEqS5nC4Ux5dcxViy/Z+FKY
5sM6eaFsRERza/+ZgAh/Oq6h5br0U+eUIzhQrONbUOCwdRLxl1a6bKb7x3PyKxXWoo9sgs4d/n3L
csIh2fr46uwWNJLJ/BZGu5l1C+R5ZkGr7mVrl/p/MTqtgciJuMHnhebaR8pxVuSuqjVnlLXDFLjQ
AfijJhw12rU34+AW6LQIrUyqPLHqIXE2QeQbq8nGacTjoM2atI4ZHtsQph1zvuWeQh4x59VyU+8K
/2fUzbuAo87HEcY5brWrI3bG8y8025NV+UFGgNH6wevN6CR48tEARjiU0Dn7I1bvfYoJR0uM2umX
XS7MiT5WG5Hj/qvhDvLhpMXojnSV/I5fClI1VmfewaHoAnco5b0kOm0g5F20GFxdwv+GM50BBj8u
Qh3S0bX8i2RBLj/ZAzQ61Xkjbz1Zs8NwmwreF7mJY3B9UmtPYyI4CU9Yam1AcXu5cqqBoi3KCamB
POeQj27vZmHEBTB39koJvfSsKnrel2mnPIFUiLEND2c8j+QHp0HZRLyOmgolucZVcs0v0e6SmXkG
xCVftQwX73zu46HM86x57BXetPjc5TsK7tUBO0bDJlcGXcEW6rug9heA1qdouwbLbpTo1qsB9Tt2
LjC1B5IYfVB+WSLv5x2igQ46zSYaeJn5sZCXihw95cWFC9C9+6rVyvP0atCuNQd8cPJ2qmVTWFi7
18p5Dy7f/Cu2++ikeFVt+WuFkUV0azkTX4hcs7buqwVi5LUKSHUTlOtBSmMx9ToZ+hGZnPcMAUN9
1ittRboMgNBhODP6aay2c0EKEjTbVQXYw5Lf4kpkPI7lSg8M/0sR9V/3/lF4nSOZWe8qx3EFEd7l
NxApYMSKNCw0h3lZN+khfd4KOvqDzx+BiiWOPCSThVGV5GDgdG6BOdKVgVB+ig/6qIOQO+pqKReB
e7gWQ9w4yAxh2DLRwozm8r/qzBThS8sy22M3puaEX4ritrUUzEPw3Hxf3GRJ5dShnWMfdxfuWPpP
rS5Gnf1WmKM9ho/BDXhaLuKcr5tG0OcF2C6yMMi3k1IcBvhTB6y4FfLt+IQoKSdoVEykKTKszMF7
rWKqvuoitqX+DHfrG49QILeV74M/MrEhkghoS4/g8oSHwmvhuzhQQ79mu59eoyrgwYpXe8UrW5jB
5vuJMa0td3hw7/vTeeT3QreUX3JSWKnqU0jE6taCuNbWsxHEKBqrzDwkRDGkcf+Z1sJRm2R+ZOno
fhsgn34crlruI7/sgHlvAoHAKdpgwREaceR62VcZ36DxY1FQAzgOdMte/SyovUOp4KcQW4m7Udls
67rqvKcYjEVPKKoC911x2l5284rrdqO/9aGVggT7wvxuSdIuQTwljA5KNASMsdhazKPV3NKExtaX
cfH7/+QZZbjaiLCojTeunx8sHav+HqJFqDcmpcUM+BKz7cd4PYiZ3ilpsLoxFv6syylYMCTbT2Pk
Ugby6xBdxAZvr+7G0KW8PRYwDG1Rpmp9Vf3dZruDZZDw1vluEAiz4/STUN0KdQs9ld6gOLGtixaV
HjbTmBlfgSarnavfhivaX1RZA6KqlxdnqW1Ra3UEtdVxaIeVmx5Osd0npwrBwi3aFAS7OM2nHKFM
w5X/hzMJKn67O91dPkxARcJ0lzT3Q/AvjpjfRlUfJL7tYF5KUDJR8I4RG2GlDb7aJ6WRHcx7JmAY
lRFkCVNTM6Hcm51MESZirwBby4pWS+GPEGExNj+MpHxLzxDxfmevb2hxhbT2EBrPqHPxyHI7rm/b
qzACf3NV/YqtDV1YZzbjdqb1UQckJyvSKQzk6rfcSg6iUc3gKHAV1s0oE+A9DkOH+XIchaxGWcpY
FfcBEorWyf4zC3qItYS942y7yiBYDqdhDScmglpW90/xqpLQLxDhG/WRPfiUsLl8iAbwFUbi40LD
ZG39eRbrdZd+kL8UfmmYqlLNm3Qrb1+CYuOgZ75dotBTLE3t2Mneoz5MhST7qT4BmRCUZrgkFbyP
buwvfwQYruRbXgrTh/LbQHPSVJPgnzKQk8bQ3JGHDGZYtvGgTblFw6GniZH3/2zRmJgOvpj0Klpl
SJPULDkiiCHRSZMBkOnv+66lcBKGdZ5P3CXBalnaShoSpWUgs9gjKbkvj5LILL54lj+zWqbs4iIK
uBufe/73I7hNkxcyZ0bt9cEb78gl6robOQQLfQ856Di2v2waWFNHfOp4OR6yyWM4bJBr7HsQqPbR
regwPuEw1gv3HSqy3L6DMoT49vfoOmngwo5hYZNlYn/I5Vv4HRJcBFwOTbAZEcv4eWbRj7JQCTD2
Y3jYZlgP2os1hvdVRVsFuH9iTPGOTUgBowuUAeQA9dFlkVRYQdAw3kuHfOXlcbs5/yOpx3bJu77b
aJpyDpnkeOZt5GFxco9sWjk70QfGubfsg7HBU/02RHuHBbtg2Hmh6dqWg6Yrwxjg66Q3Auj3oS9i
hOeD51Eox4hmS+fofUU++4JK7hwmrzG8N8Uwqo4qyCfOtUyciQZGak5i1xSIjwY0iD/zHg9Z/ZEj
BVS8pWp2pxxBg5Yv2YGkK6z1eJzNdi7eD5SUyMHXmn/eWuvWY9etirivwRXgw2+K70Md+DNx7RB/
ZIzd+9BGGCckzTeWhazKF5D6wVV6NbrMZBWz18PpqwzW0ndMdD36PVHjFAET4VwP/NMjCmlxB3UN
mlF8mrpvxwlfloxgnPJvjlhzGwQRkU00gPNcI/AhJiN7bgRIy8CjAMofD6DUBvyJjbcjHRaRxpuH
XDJh+h+lUSFidWYBFExtHLoHTLpzO2U3UL7aK903LZvngVJc3Hm1BrsgGGZDg2QwXdkUImLCYC9X
lBOgOzqUiO4DvOCRKUaPoU5jSoucikGvSBakfPSnMv5jXR1mPiwb2F7p4ioYPBFYAUoOCK1bHVzD
DGLNUBxxRVz4oVbC0maOAv7WM3FMJrJAzhbWtcxOixT54U1f1Pl6emvDIy/iWAeZVc3InrV1KdJl
K8oFtztxEs8XRsbRde+PS/P2jfO0dMcoaNhTrX/NZ+/hfwPJck3Tjsjje5R+0e/7lXSgtO60+Sr/
eGEDl37Jq7rKvyggeZt6/hw9UjzWtDMxPyezROz0AVVtg9ugFU2AThgWht7jaoSHm7T15wefACTT
2uyufSsTgdWxnw5fCu/GAMA2wAtPt2ocA0186LVTTW7+bhizxvmGeQ8SWvAED71HNCGmFzu8vq9o
QnDMtKdK62iGp5MKaA81IKpxhkyreQQRy/p7FbIKSOQWHbcOkIJSbWSm3Pup4xHjw3VfkSuuyZtV
LA6gApgmp/d5+9m2u+O6gULQJJRShoMj8RssXhzOecInKv+Revppp5GH2JW4IRbtKMrT9vOJCYZn
f/hFpQyoFxxKG6pGab77yyF7wzUqTOSyztQwBvzUakSqK3ZGzLAQCSShe86KIwK692JwRgF1tOrJ
ePgsrRP2N58ME4MnTY0WY6AwsuuQBkQugHYrXDHDFu5svp6Avl4sYmO6UFvHJf3zbDz343Ynmd2T
brmSxLJheuKwo+47Utge59YlnM7bk3C4VSXeEHsXQ2cEJlTnq+JRX7kpvM2FU91eGn9YMaFB7+cJ
RGRt6kD/PYD0qj9c4l1S5eCe4OB8SVdojmAyIdUfSVrV+KB4yU9Pm5thT5yzi/BsIfVqPrvOa5VA
kFrrRMMeq+y+9qxj/ZyrDFkpLHPzddpqnl+UdBJcIl7dauCZEhR9bjOxYOud8cTqolKAFEs+4iVx
qjwJtReg5VKbgqmk9XRTIM/UkM6aeVfRNDJvGq/yJlNjxio/lOeDu1bpgDffhqQXhMiTvUNBPA7Y
aPaOcbtT1L0pFzGVGf8+MCW+Nad7ajBsjU4ntJ3N/ThcWC6j3A9nYOy3XhZ7fMzfqsO+ksZ7uvKr
9mpeseKWV0u8HhS3hHVeToO9D+kQ8QSlGPSk7MKWrhq8SVng/z3UScBrBVxi5pwlktBLftynytnC
Ggj+gp32mcAbZLFEPALfGBXu9xzvtHmr0t2QjFDE38szjzck5LrcvF67W9EVU7z7B8njLij/ay2c
urQ9PEg/JpB+S9QWA3W8hM8fq9wULUots7Lzd3sdPSkietk7OifYmJ6N+w3xVcbtb22K13Zv1yqM
amkKw9bDEWf8pjhBxVu5dTWH7alWFwxxTEv05Eqa+IPVxoN3G4z+FPXAorptjVrngo39DpYo0Sp7
Mam0sCSrxFBOKKTdXNSm04MRGjfOkCTmgtNG5WYsSA6RqBDfD5jD3tzFHUzaAkl45Z9w/a6zmDeJ
Zzdtl80GmEyUZ15A07lM0Y/bEX49ZI62DynJ8f3HZYdlOjSDWRUZ+xCyih6Va6avRnhr8DD9n8/y
4DUcWYvUN/fu7kmmRAAr2EvGula0B5GZiBUtWlCEI4ZV5/bOga9bmRVH6xsaYVIM2kP1lmo7EcWq
JQ7VcpjFsQxvIgWXk3ziM1gMwUWY+vKH2YA1Io3a4VTAuB3oCvLXDKjVqJkBjX8pcAjehdgMy09+
VNZpP2vcYFtRe0gzDASlEnskz6qukN3kT33GSI6nLjtaW+2jQVTSOOrZ865J90cixp7I3qRq/hbs
aJAjz8yyjj3rjCZmyiL/Bnl82ug2hc+qniNof2qVyTNbbKV7bzpYZfGbCEgxVLs6aLs8J6htVa+Y
I5KEHRMUZKNYjZU6b4xb+a8mZEP6hjJ8dtvD76bGvwEYl2qFx4/93aTtMuqfZiMeIsxol8IBprOc
DcedXdETKkx9vLo2uGQZG0sOdsjN/iD8wSMkJ3BZ+CKi9wjwakwcb82zCZWLvGDTfBQlEdIGnGJm
NV8pZ5lDuQ1abtP6McmdfPj0Ll5egbFY3JDKQ7KYaIp7WejphculbY0cktgkN1AT7qM7W9AtMIe5
im426Xza8r4E5b0QDeLlTHXhEHvXNMjFuOKfjqkXM/ttKJvDaOKXu4NVUO1/vFNdrAKJ/AoWLBAw
q+eW8iVg2dZJyULFScQ+esJh+sqMmPNvEnhd07+VYFCPRxHpsTtz33+4ZS+/f55DMp2//2PRBdat
ziZfSiY2ngbeR0qKWLYsjxI/GV3TpvlJaKcuvjJQWuulswlNBtYPeV20qYVbseddh6xquuLSpVOH
K7VMjR8uIDMlah+ztrvrBdF+wEtMsGIm8D5kCX9mRsCiiKpZDwa/TqpdoD55ycnFMxP9kxwPwEx7
z6OVd0BMK1iaalBuFlPQtdtnbADZybG2mItbbC2T5TiSS1lkBVkIJPOuSMPvpduQm+Vv73Bd5FuY
YYqUKA+A+ggexB38lof2l4VhYJUgleAQfW0I9yaqJLKr78b5YXW3RiigAmkAHx0gtqkjefAWmhAV
NmpZJP2ijqMyA2SKKv+L42SgFHVnoTaLF6QLLLJ/CSJu85PxgdavmD+PJw19PzS/AE1cXRrx6mgH
ID0dcBkLrCpjoxFF5urNmC3vOv6Pyp/gA6iNcKT8jRD1kNFMt8eERUFgIkoqCn1s1F39g1qA8B2W
K/+m+zAVIgQ/Wu44R3VFsdwvb0fIgPMcL1loQGxsDtzk0juLurmXp71LmZSIXDno/5363iQeXj9p
gb1iYdaG1SKfF4kZMkBqAlm8Psj68DS38IDSo6hEHc/ho6jL+pi48EdUZXeLKXJm2N4Fq9WTghMP
iXYOjAu6xwEJiHszL42rV+jqml72fyzbMJa+bJgJPLDP8IjKlzWpe/TONhaqOOW+r1L1VaVMbtqZ
XPlga06gzwitTVHW0ToT/pNpUIkTyL3TCPmaVqwCTzXwMStIzyd2TrDMycgR1+ofZhWeQDjNk3Uq
xRqXLWQFHV0Zyk1pYcbz+MYK2o+uA4siiuRtRQC0pHNsYIkk2LThwV5cPKVz5ip1Uw46S5H3FfLy
jlkOXtLVm6mxCFxcwxU9f5RLCOs1BdaiokeT6XfX81aKnJFqGKKlz0uDiDPowmU2AA5aCQQaa+5/
X9veAqHjDUOh67O+4P/LHN14HvWCr1z2W+Iq5v33uiBFSuJjRCSrDtkNyB7fFmEpzJgEZ6PQKXzQ
aX3NSizdxPYjc96OQ+YmWQpUatGpze1Gh1K17v5GHpeOOK+jn1uDVLFi/OWjO9eFD3d3ngP9jHj4
RkjjSM35B1jniclxfcDqfUnSOrfbGuNPHtX0sI0k+kSn9gSbCg9KItowKRWFvDvLOHFSgk59ucd/
AdFuxnaT0DqKPD6AP8lIqBsCOCNYY9x0+w76qu6B23SuzFdPT1WrA1E2kBAILiugllzGMSRbz//9
8MBe9Zy/g2uJh/ygqQmSshPuw15oMAMPqLRZwV3F2H/UCzE/YXufyuG7nEODqXTuFKGFvaAi+pyb
rW7kYU7d11KBpPn9YpnfCecJsOzrjzwm2U2uRptTc0SfoUdKrGyhLxPk+1qIpS0EHQdm8l2CD04C
d1jfKiG6g3ISon4kTYJiE/WAo4EaRFsPS00etMLNWp79zkJO6xVJFcuLoMEW4GJdXodk4m79YUv7
fcx+WqJBCVHxIVbsB7mwk3DLMWjQWeYYd+TRmOgNZiyFKurvavkW/pC9zw70hfvjx+70tuBZm5gM
dSWI8HqpPjA6PckykmwU1nNthAa6S+oseqF198GPwUYu9p9vgHEUfM0rMjO5X1tu4kCYJuysrzvV
HAMnVxu2fbLMdt/y+Tur+8ij9/QDcwL/S51kRE0rfSSjyin3PHjSl7eA+Q3Vc+quBMemakunaXvv
Oagd0qEvSbUWJ8T/Px6OYBtKRvzP8LWmLB5xTSkJ/PfqJvJUkmiAGL6cxUD4UmGV3tJIUdYvXNLE
82r/htElYxNlSNay17Dadtlg9gUka98XCpAxymN5Bv6VHIHwOUgHX9d68akiYCSyKWxiqHlr4jYc
gvxXRaJDPIrL0np3WZwaUFTQvRceB1atdAy9C8SGihYumrLxj3AfT8ngo4rfGN6effjQ37iXMT8b
pb2PFQ1ZVBA1KMBw2xchRLgGFAvhp8kM7qd7MC/SgbNCdJ1PeS53wrf6hyPi4SPWIncw6MesPlPv
5cg3csL+l4VNUENkV6sYLVFGkvxYuBMYUnqdj6X2igSCUdZ0BylT0j6RdOhxfjrJryacSN/f9gOX
iiAgdYfnpsuSDRyJRuDK+8aq8nW9o1h0adAZYaUTOvOnF0a8CWqyIawjFS9os31zaxtHqrf6Us5c
DeflMH3LaoVLKH3kI9z0rMWVFB6VSwE8evt146GvrMd4apHZxXVlsLohJMzgp/hD95wnDogJp/+3
xSddppKvhTsH88ONjF7CTrlqyLUPRvf2UiRT0veFmsbUMVC0yYNkfUMHp/0jFvLyHNnu7A08whvw
4izs3I9QY2j+Clh1mw5w9OELPCYfALB0dg3Ao+1cXBoYDyPHu9Z8RC/m0GYaPv7bHypQ73FAMH+M
YAn3kY5zHdKzdv+RXPyjG8HPP4/FAuG1NI2FrK8/T2xFE92b0N1fhzzNmjx1DPqRKLnVN2+gNq5Z
ahvyxA2fMHGhpcus9WiGqEYxpzOt1jla64CwhGfvZ0W/oHGy/WW1CvA4o61g7uDF267yK5iaBh7d
Vx/sM9iiaOTSvFFio1BRNP5uONLVCZbnl8+TUXCl478lta/Xcif8O2ry0NnknvBuIUTrnqsV9I47
KTuxQuvQr891r0oSGY6YUmIvk/Oy6HHZzNSMNvreX894Zj96be1mjLkfv7tir4wm/kYwxFkFq1NS
Q9mCF20m4gkaw+X+2dRYf4ihJ8lvlaGTPkH+SFaBO1acixUGHEG2x+sd39aN7IybekR5jKj01H/J
8G0Dd0jxa+X3ka8gl1tOtic0SK3s+09lEYx+XBArHcEKjeag4xy7LFMWsg5lR6rGzAt+/N4ZaI4p
qzLQ2O0GlcTKQ0RUB6JVuWvA/qd9GVCP7l/AKmt+IephHcaSPuldkkIJuLJWHq95aghJ+FNiX7cK
6WlDHU/kxGT2azdv29GIg4FqGE981x62pFRC6J93C+XaZVGRbIObCCZnEUAdnPQhqxnSfof/aZXo
WqnCpukBCSJNPvL2VztT98FkFZAAIVt1SXYsQLainsT5Pg8CyfDzwe72AP8aaAgntriEA5Yr5Ffn
lzaYTJT7eZcVdPVh+0yDbDTrbtpEXLp05WwlU35veV7s2rPHqxelgZRmV1kLo7nYuO2/APO2bgMp
U/KIrEpEO2aZy7Po0XfGib2OHwPArUqE8R649UIlQKIuzhlHwlRKBqLJoOIialIdQuGu0I6fkCsH
sgVohQfNx4ZXOOo9P+dr2g57PU1uHeBniqedo58Ps2iNlam9O8+04WuuKTQp2Q4ILUyBEWY3Smfj
mBq1bpD9LXKx0bFY/GEAHoA2j0/FrIE9wM4Yzg+m/T5KZHRuKO8xLM4XGCKLDNdOqBdCeiXyH5rh
YrihWJuYX1/j+CbZ7UqMQXnWPXhlXUnAT1OI06stXyQMRjSlRb9ZtfqzZ9lQkXa+JCMyFKiGywg0
seV7P//FsF+LgxtAwhHn47+1MPGRy9C5V16Bh27Ly/B4ZJ5k8BX2SiDnGsZ9RO/LUfl7qtuu40yH
lNvB8qz8MzhekFNxk0iDRQma7e9gfBvMY9hAKdNKrx2qeYfP208Ktjm9scer9i+LoZL4PKEIsOky
EWxmHKJyH2vLxyJhNwD9TcRaZO4Eb73EtAydhAptHts/VYAJX+eHjlwucr/Y57/iS5sCDyoMW5eA
ON44o9d5PnR+na7St7iIXBeWXtAN65b9hSA4wNe0qMwCc2x+FxbW6GEcg9qfEvAilxc8T5+/lzNe
cu51b2b0AquX74WueHnUFqZ0J/xzmzWGYVBF2Wy26kUU4jJhv4mZOFkiHrK6Aj5G+mIm3j03XTOH
EsH5SGYZMrpgGqGNR5Fh7if+MSYV/2sB+2aFhGci0ek9MbD1/f4uYBfCX3E1/4V6dOnwgthsvh2m
ASxeyMwbBVen/ihWDL6jLYb1KcqSOLAS5rzMc0e4/B3Z0TUu+TftKfvK8vzfZczvab6Er4Q4JnZK
2Hq+ayUEau9jd6FK9Y680khsVOmEf91ke73VXr17z/RzCNv8doTbw1pPCwB7O+qaLqK0f8EHqyOd
MEIT+ndkNYgMEp3t2hQHQw+I+N1RB4VEh0pP3rUgzg5tdAm8HezcBdLQHpfozVbALQ4zobzdCX47
0hupj14VSJx4fUUU7GnGOXt/kZn2vw9kGDRf7NMCSLn+K9yU5tWyF/ZaLYQHBQZjPUxrF7HAdqgF
RlSLd20oUKOkpXU/vsrZKrWOYm+duy0PegotumUQVnfog/jBbpLxTv5XO4g3UmjCP+ZlSsvEyvgU
8Q+rXBYBW2be3xlaNuoqBLFosD1cqtz4vF/U0MEGBChYxO0Dol/0AwcV/JmGk6bWEV+laJCV+4np
Riomd3b8+cbsJvR2YJprX2pT7EKsbMO1FDSMEsKHtb80UBgBY54glTh2GmTuUuZBDsRN5z/V0j8+
gImASEVmljHgv7t/Kk2Mj3MJr0ucn5i+7g7SIAYsxKy9lfwdyZIz1ibD8HsP1WkHKsXQiHiW9u+9
aH/1tCVsQBlseadRHWuXMnHoe5HWxSdC2F9dEtqQOa4smnEaXV663/HF4uAIXwJMwOVcnjHhiuqf
T5yqVvNgnTBPMDOMyA47Snx3aJ+bPlUAbelR267RRo2lMwC6K8lb45eV729RhbvISiQgdz5ZmfLW
TlDRv8ZOxVV/Um9hD+JA+pkmUB+nZIcRvnoeckaxvtG2ZXkniIhYU/T8mDeQVwuWYZH3ZcCTlJ+S
iBXaEwpKaGLu/VAFt6u9/oQq0ofM4G3ZABrsKXMCnXRnhYGkr8wS9YI90ZL5eRg/QFRvPlA6q4ZB
+/zOtV5HJujs1bpSajHxvri62zawdFKbXifHRTtlx6vckmqa4uM0Widr9CtHRTNVatDPJS69Mypc
BzKZdSzSK/+OfsMPwsIe4ivgH/CxM9HwLjcVzgWXTOw5Edw2inMS1bAvP4onMQ2wizY8KqHaGpnv
OgH4dzResPywmAikNtTkAF0hYP1MR4ymG0uhJkAh9/R7dvrmVZNBDLA5GRp+YYVgnbVIlh8r5UdH
k1K/FReV0gWgxayzudv2nEuuL0zX0f/lYJaMigKIn36HGkeIzADKRX60DJfL6EyNNVEkpagBHXuL
9Df12r2Riwcqb4LFuUkP4CWo5cE30nlP+ME502ydHuNw15JCayXLRrHbq1oI152TkSOJlogubgrP
qKDSrX+78uBOvghXdqtuyz5/J8YprvCvBY/ey5YUp9okNeHc85kwIUPA6x3lJirbKM/zFFsevSkF
84yDToYOHkcEZ0tjbDkthcXuXW++3EEaWKIcG86qOOPOadVEgPdnXSjyHeoyqrQ/vYBjhqBcL1qr
sCGPfumDMjuix1ze//wq2BpXJdsuLDhxyIPKQSxjp3FvD5MkCP5GK7wd1uRsJzUFttjNGcP8H9Y9
ciPDNFjTt45aEk0pb1rnkz1f+7jQQ+cN8Hmc5aJ7AQ4oH3KXcRSnYqHlpIbBLtKY1lDXeL57p0WI
UpVIlRXeRM7rY9A1VvZXq7KjyS3Q6afKsBZwwJusVHWnHZ+rf+gaxaqPvuR0J5CEDagNX71N1B0V
G+6WwSHrpfZSdY8+kakVulMI+Cm+vjkNq9kLCTX0rsY+tiu73llk/m3fzKqg67tjuqndyFQo+qxT
w9E+nBYekEraoTBOWJ8rH5T3cwAlrshAB678OyiP6ZdkIEqBDRBKAI+3QeJdnYROiS23aCceY2rF
Puw/bX+2zSOf0rxxFl4Yr5VkUsbgJMzkpzKBAXVug3eHG5VAVtQ3rRqmOV9s3qdDhO9r3DlTGCVv
QaZVQ3SnEzE2WHTzSIKcj8w2zkUOhOAS68gHYz/Gqysp17jL6ljhr9XnwRACx2y5xJ1QbYGf3uRe
hpTrX+VIsSYD1lXUXiUEnZ/RE0YOMS1QNY3/iiLK5qpN4whEZXEOGe6kT7KEbF7XnyztMmEY8G6S
7dfMAAqRFujADx8ZzTKxbQGzAhCLtduuBFK+5KIzlAes9qjPrteHFrL8P73Kzen5vJZDQcNRTtDQ
5R5wkyJCY3i1fCE689bbf7FW7bF1HvruoXRHereq6Ctot8HksqnZeIdQGWT9I6KLX+em2IvW+xsS
uHrXP8L/oDws0GQDnmGRWy7CnMb1tbIiDK4VfAk6Q0oUMU9QbhJOBulpdSRfbuF2lem+NBumYrbU
6c8rZ5rO3kt9bi4FX/Ke6/7xYaZp8izFASEV5yVYmDp/9eTbAclLS1vNh6YGZiAfAlMCPDyT15tn
3y/BT06kwoV3ivm/1e9gbepyyN+dpNMTxiK5SWFPwzbDBe35y2+N7cPSElg4EcsA3gKqWkQMTxny
nAjk2Nz78CroIt8VBWzOEDFCgQbcCJQ/oK2ilyjgnqT8dfrKOHvIPrEUaB7Ljkx4yzEm7q2DjyXe
2olBxwCEHZXtcE/JeklkYLeJxn/q8aUcIqxIb9nD+Cn7yJfmSVgoi8hT3ZUJ+k4UX0BZLfHU1sOP
dU13xX90DCVCRoKDN1G6e0sM+fRucfMWwglB1z9qy423wrL5CkAOwXLOoxTUbWPdkNydWwnRHMtP
VHSdQdd5cINzelKWz2tMJt7zLQuli69xjnWa6zj9RTGMTMOYGj03yC7D1bAP2bKgGl9a5H9MB8zC
HAMuF2s2iptWyC/q0RY6kT47JAdSI0XEonJ8RIv1p5NXUqIiFhsCh+1SO+T5uxRJANCY9Xx3OEpU
MW+KdFeXtJp2yE1mLlKjOP6ZMzrfG3awTvp/JCPhp1PM2XsTJKRRLRwJEz3LBD32H7yni9SSnWje
SshDv1/B2D0a7rkTZ9m1XExbUcOgvUFSocSqwZ2gIquXuN1KG0evy1cj6E2WzsJrixR0Hu/T7XSs
Z19nPbAzxWs+hvifKwMtGyRv6ja2Fj6agHfSwPLTDQpgBlenoiemuJiseLgXHu8QlBHErRiHZ3h0
86NvWb/gQXG5HmTRFAN/VR0gybKfh3mZ+PCexzSRaSSovY0pkvORuYBytL366CCrejcFJQ+dLjQP
0H7F7t+h7fQ3vij4z1ZK0igephki2KADJSuH26lGIaaS/x+VxtIRJsWo+SbSmYFY+7QSI3C2vysd
vLL+xygZ4fB5/y5/LTB1aAes5MDgyi4xnb5Ln4VK95Y8G6RCZoWeEJxzb0P9/GENCAHCBulw3rEp
GRQZk1JieZh4ht0fFKCP1OuJqeaObtRs7hBS4k1GX4CVXK3W75L3Eh6EvxStoiCzWoRGuZljwccr
oSUEIJTfqV5bVv0Se2Vtd1JjIkyvG/Yj6EMeS98Ukc4+gu6/nlHGubKbtgG3P+jK/CpDSQMhGKk1
pjNK1zhY09iWczX5WIEpf268wW8E3XrqhLPBdtw3LmyhI4mAbDCM+p8XmS8tSCft6y1h5965rThk
Xt8g+Srq8uWrbwzdYw1XYfnMySR+ctKMKvqCCA5G+CfzC+YE1Hvdu5/FFK2sVP/f9dIWw9wfKtcw
bkXHGqdTOuzBO3FbZ3uQ5OQaXxsIKqGHfc5acyEuNz0JwfslAOhFaIlVug9zC/3kTuiHlh9Wi5VG
yZsr6lMrlEgEWWsbs6Nki0JOGEcA/Ch8T0aU73BOs3ZfRRxN7A2A/JQs0OjF2gL5MtcaHu1K1dt9
7CUPEOnJzyG4a44T8fmIAAofmlxryaMiynqylla+TAFzXEuzY1APbfkcu2+HCL68uG8or97aH5L6
el5s9aSqxnvov8zJ7zPg/L6LsA1P7yk/ZttnXNezc3WJvf3jQLukkaN92ab0ygPxiCPuSFV2p0Hy
dFE/buf/sGDvqmqEFohnp+LO1UZRtaX625KptPCMlRDt0K11WIrY/ItxCPO/n0pZsUGQ/eAFwlqa
cgrUdOuLPxvq3T5Zh3+8nt04fl1bSgOAGx2xW/JpLxrfGb3nUYb06IKMWijF6NEnizEE/I7D7dzN
hgf9OddkL74HzLZ7elqIHidcgL5SQzOG3SWV006UCwH1G0gi3/v2ZpOdytFw5/f8R9osJvsSi8Rh
wkpoSGXLWfwNlQrQZl5GEzqRO30VHwREkBW9MPo9mAE3zU42VH2hEqyHdeWtmuEekwklUdMFmCkE
DR0tFu/jAE/kdPxJ5fZPQ6ZoZL8g5EREuMqwvw8rI/KK2cXaVRdH/ywRhwuksqZA6qj+u0Jeq4kw
f/TvL3IIf5r+oJhB1+D9+b3r04j0/62b6i0oxm37H7Bmfn6RlPMqG0YFPGClfKn4XOqPEwoZgBWG
5hqmqD2FSHTIBui1742aMiIUECLPtc1b8udd1m+fBwuHoxwmnOTvGiDRtEwOEurL/AIKm7h+0Ibx
wxxFybLSCl1Udc+iEechcMN9lh97/KUgvTpx4o8ivC/HGci0CbBrWUpDVrgMJxVBNdCD1xHwmEvT
4fRFNkhNKCBtBwSKmbpgbGJ2F1oeUCojAtGjm6/vL3F5hnfTTKCveQ1XjpfaBvzCEGG6qpbmjBBI
B8+Z7pmNmPDx4H0CNgu1FYM8ErK+4+Dg8ASudgEQ7fdqP7uqhhzY64ePbcnBAO3y9anrPal87HwL
aYSh77qTFpJMFUriy2MEbamNqkBNa4kBPAYRhAk1dR/g6di6y4BkFsLoHvE0YbKFJtyfhmH79qg0
fH8q33OWSHztKWcVjmiqatRwy3i+ZfvBoz09lsRIxIjPBdvMrlPgAIm2VodWEZLCYUmjwDNJYGdK
0MgTOqnzClHZaEhaBdEh/oWN6r4zEiqe+bw4tg6njRIesrQGaXhso4W+7LTeC8wdToS7EhtK2u3P
4iX5XsvBB2msxHLW22H5NGahPyhf78p5bLABl+vqZh9EoDe/IGEIAY8qk4eHq2aCkDb4y6CGRxah
SThPDFL3u2u6PYhS17ZMU0FFFMCeBKZHC7K5hRSlop7Z0wRsps0MwhCD4l6vCvFg1Inn+bQneVzd
oZLneYsbCbvNnmUtYCmv1G7CeThnkj0U4HPEcGPKegrmKOyy4zyeWsGPXmu2mGCnRkRFgkitHP5U
icC0wvEMvtpO7pShx/Qb+nmLGABXqTDrrIQorO7ATZhW1PH182aJz4JVNQOgGjrkc7KayzVjoeAQ
dZmnWt9LSCPxiuOM/kHsXaHxJfTV9i+8fdDyJAmUnbp4mpBe0t4flU7IMYmVa6G2/FGQ6kibjwg7
q2kYJSFwu2RMgvkKMymipgA4dS6nwTh3ct8zS50XjQwBcuDstGqIRvd+mkPI8R4gDjW9Lv5MaEHk
dbGSOBZSiSYPQAkLjn7rERweITJgO/HH5ZougKo9v3cB2cInNHh+OjW7vlLZMI0FwIVISI1QcZeX
SXkvfticxPsbWFbDWTsqwYh05c1uuhfaCXO8otwmaBsnpIPeGbCWcdt8oEKzarTIdiAS6QbBM4AL
64qBiQVxTqbfOQbvbp9CUu26quxTE1chE/By44LXdrBx0gwQi6/Zg+py+QHSNf5qHAPREC8N/In8
lop8zD/xT4Y5mAflDRx7ztT4wxkg9oxv77fA+AB1I+evl39YwE7nsfdbR77nS6HYFPqmRM2HCAHP
PajvZcUK8WbBxu8lcg2VvO8aBUDkfPMV+Fsu+tQ8tsgqbFNKjl0geBwcs4PYxTznkb/aFgptSjqy
55v1Y16XgmBGARSvdSeEAh4xGgwWS4vbOcf3ZK33j9nAigpi7Ouv+tySbP2+K0CyzePYUgVFtMaw
AQU+2IjSTiOIrRSr+DQN5Uzayf0mf3YJ+woU4Hu0QowhvN4ZhopstQpJTDV23Rl9KPncUd0dHY2K
FXSFGVPEjt/zxvmFu9fm0dATwpKPDDmnAXZwPgZcLaNsgiSKXL23NUKkcovzF4cZIxvGkVKRaOD7
qPMSO8Tup+fi74Ecs2rRCP1L0CbJGjryqU2jOev+IeXHt84LFhwcU4hDYOW7Pj8zNSH5nR5mpbeW
KNtVrjqJYgDGZausAAxLpMMm08MdogF9wf8NO/2vUgph2HTC5wZ1acQ1SXKL/9mpcn2kR7SuSd5R
ymVTaxV9+0V/+gVjd8xl5mLxBoK/3LnpI/eBpN0iw2fsdqub3GnR7J++yBtOhf9s7rBiA5T80G6L
UnoAmfV7VWOEGQmp7q2yEC3XcPTLJk/s1fQBR/AKu/dljEf9LrFus1SYumdtc2NcUcJmIAUkIzfB
qic/iwWtZl3VOcAaqLixZzlRLJXqnrMXE+ORpX2rNSIJSqdsiONb0k2dNLS/6vn+1uAg4aVCnUL6
0ojPJbum2CnnEwc6bicUuXLFxVyRjSlxZ92SnvSvZGwx5V5MPuhjvWCOvNCFANrdlT4LwbdihxM/
q7JaSRTAbJPuevlF6MVMI7FAlmmC2BWmmlr2OYAecIQ8K5GNCvkUMiYs1eMJBc8ex4ur7S+yWswH
o9cWq27p/XMXN28gEYh31cs1gTx2dzPXnR5U8uW1hRYs+imZ4gz/OEeixtntuqfcxk2ugCWhZRgG
TNmvDIz8NQkchCfGl9YXJlvjh+fv7jiOuhYBol1vNlymwLgol38bD43B+ODuTmOOavmSgGctPU4z
6pUCXgk71fHSNGm5tW7bj/jarWv1ShK/SlR7UwaMBcxqzDiXUt0B9ZzOn68jDpwXUle/jlxcR+x5
0x8mIcZowxD8f+oTDdzCSngH6JpXz6e1wGsq7Bj5TmwX2HDcOoMPYB1f7IRqxwSp/zaZzOCf+Z8d
BiEQusjQt3uwwGhiEZJsSsQlGyoBnMUnfSD3C7vEVi/m/tWPH74FTyny/pnzl4SU4KwBFGd8x+az
egQeNV2a6cF92+aj9Or4ZTdeWC2ZNSlZKp2+x9E7NoZ+joI7+BP5ZxO+PHz5GBJjoNzH7oZjkVvl
d6Syxf1nV68WD2X/MzUNc+krZnX2Rv90WRoed9bqN+CXlOcD49RY7rX3x5g38x2/VIHTqviLw6Z6
tXqd/mP9zahIXruDlkpRu2MebA0c1izaDjgjYJhsQ0C4HNQG9pHk2fMoIr3pxpC+ZSEBihMvcB8r
32HRELet3mEyNbfzsChGlfSbDhHZhjq9MKLdjRSUy/8TVU7fM592f98XRde1bu7guEHrmJDPip6+
uKJnlU9uYUe5XuLTixZwKNWa7f1E9V+WdLyz338dKgMw7MIwC4slrP7DawitrAijg+SCqjXY+o4s
v9YQmV6iZ/pDV7ts5oYEFRyqx8IcQk4YXTZBzhtc+zND5/nQ2iTjrtNNEW9jASiR3uN9T0imKza3
sbJcbhBRMgRiM1eEs4jgY8z6TZ4Js8oaj1GWhuwrBrERanJOLxv+XQmmFifBmKChNxxPuDPWPa9v
oXZbqDGysgJjnGve97w5pevdDDV/Nsc3NnK2ChwTeUT1DCfYw7qXxldE7SwSKGhY8dWWY8YKScyn
BtOSlQCwRKPSJw2TOZjoB0/DCTZo9s/HRCjXbl6km93uzcKXrJrmwoic0yfMe7IYm5tYc3H4wcwd
w3moQFoPoWY6pSofNZqJTzX0qythc+vVgHHb6zjibXbO+gAQSRDuSdX8tgdBcaUxgH55xTEp1lXh
RcBFKNMYh8pGlojdpl7y6Xl6sasaG4l9KqQda5omlYZWgxShof798AApXhAVi8h86bLFX4m4jhmW
CF6j1whV0WQVaB1N0tr40Z4uIqh10blXjW4Wm5kx6wzQ+I1IhxzlvPMAXTy2tk1MgfYyDNAHgN3+
72aU/XGAJTtAQxusFlxbvhkw+diveF8mpDTUxasedhst34cTB4ghCJl4/xWxA7RaxiRjMVWB3aDY
YHW8xsfbTCNIawjTsCWDv3tWCwcaOGF33PSk6c5zYMzg++87pl5bNN4rTrLdrdFzxVumu4+oUOrt
HJcVkIBvXv5J2eB8vNzaip3FR3VdtRG68uhjUkXw/FznOGzQt5M2kO69RiAs3FUCa2YXtR4MRQsC
UL6cL8DmlCTFaNS869aruOgmUJ13smM45X0ENdYabfbagRoATF64NaHsaV3iDlbPZZMlmaHxauqe
nyZ29IIyTS7PAZScvg2Jer44emfyTgrajk1grZsOoYu6d47vmLAdLHRcHrkgnynO4sEzJPoDTdWF
vGyukXYQcHEFYnpOLe8QwDLEL4gDLtluShtMVlNoXLXHoQ7ncVRPmN6GUHBM4afS2y7GQHA9SbOa
R+FcD5vi3SAw0owupjC0kS2Y68bwDP7JtSxpfzuF5KiFM1R17VwGHX5Zq/D/a+IahqkXMRBhH0fr
xR/vr8k5RPTUCDhemHxa1038T0LPeu9oByCOpG2gTrGaH/Pti/P8hHTvdAofEZ+R0bo+r4kCW5Uq
tjZujB1kvZ+GHIx71L3m3UcaXLurvpuHYI4mVuDv6NCDKsfLWnvB5yKKjp+L4+3BZFYkYmkXXv4N
XzXhC9/ME3uQYmNSku5fQYGBqW0oCMFR4ygDxQ8QVNKYm7X1oKr7NkvWkJF3kTdnd/AKabUlz/S1
5c4caIFPb2bMUsL+H1bPkQf2bkUaLPqsPha8DsFizZfDSoWkzgCkSNrYa5ismAqFhOL0B6Wmzuqm
9uGjIVHU2LzoXUHRhGO+uvWIQcUQZLYtPYyaFb1ziqKzMBRK+Xm0/x3wovghpBlUggenyJLsj9Ls
8djGAiswoPLmp44aD830pmmubuKWNqPss0s3oGcNrd10cicZIRaT93kjz9UKB/cz+n+YIumP5gLX
egGRTFVpUJgQU5Gby9QWEhJuzmpaUr7JvMWLsAqr4wV34HMMui4fowym9voXUEc1/EUOp/LpyuGi
K0WgmTOMgZxIqifrjSF4Y8D1UWTqDZFtuH93AamqSV9dpccHrh22TBO0g1xWgMbze/OuXEVXxCjV
QeSmfbW4Qnpw++kSGGHttnA5T1Wplmduyw6luEiismGV5ah1OtbZj38R7bv2FTHNSCOeBa7qcHPd
COiZjmznzeaEbyHA7PGvwOvK0a2fY/bqPBPBO3ChKknjv1dP0guu3x+0SrRyt5dP+L231Yqfhbs8
2gNwlUtqRj0iAAuPBG0FfLuHiuJ9sjwBguzCIJtnyjSiLJy3GnP/7u8l48Pm8Y6EVGioglaT+bTK
N3r6uR+qbfmnBeAofUALu+Va5oBTZpI5iv0IGBSGEYJ9WZ9kmMpdDwB3w671qcGie30CPgmEwE+O
CU2vDO607FlO7EspeTye1rMqUf5X+R/r2XwSTXdYLcqRU1ViioGyq61EH2hZHFZ8YW243XfgeblU
WtQhATc/X0IRK1jJdJBsR0q6chDCt8lFZxZ8/Btlx5c/oNxL93f4mA5/xMbnB0aez4/shlHFUzIz
4o5dFACsEtdkKN3rygGj0iI21PtV7dsUSK6Q53oRZB+7iCDO61/3lKdxw6XbQjfbLJCu2ApUkMF4
hkAXmuQqT8+JE46LTiQs2e6k/ESC9AMwyIGwquVyRBwN6PTHCN+UXTzoMBrECUZQec1bCAWkYiTa
MlNC/fmUfUnDPQG8eRq4pcnn3cMFbTT5yLAx+We4vK7oZTLWOcFMBh12901KxXZUhmqw+WnNfD3y
LUCqUrSvjhMkcLCH7ScOa1KmRLeO5I6toAAnoqmGbaLuffmv66FjtQ6mCtUUvZeJ+GPIg3/ghG6v
I+p3MU3AObTWuGElaKaiFwQv+CBAmYgIKCkXhH3Nxo7G4WCpIhNao5oOz/NxmEwPahzlzWKm7XqA
HuGCM290zZfToxCDGR7iEdk0WEanDzkrqaKn9uYIvee3U25N0wLKNFXf5LLikzfCjJ577wPkFwug
WxHIZOohdD86BbklNVvNj42YNLd3isxlSbxAEzcT807Xng1U6GyQmEHnH3ZBtADHH2fvFRljDUvw
Ffewi9I+5q/j348LSggMrAHcWN/r20hEYAIl6iDegg+02wOK//wyo3v9Fd1oQ2ROV7Td8GhE/yIv
zCmloyHePJVNLymQUeumxZz8s3GSijzqmgsxrM7mScWI/lULKqEhWsQshp62rzatM8xowBlPc6tR
+0r4kOo5tsL76AGAU2CJaRkijPCfW16Uoni74uY8+ihoTZVAKCojIaYN66B0FgPFe+6/gT8vRyIo
/xQHYW1e/hF7MkrIqNAP7OPTOAm3uWQ/igeeMxmy4BLVOtX5fM/RXucNmHSb5IlkMH0jJWTKboM9
SSX9vrJiygCl/Y2BzU+b5Y1sHwNWAkZA8Y+OD+7zTqeXeNsxTckB1MAcURQZl2onl7NO51BGDtp/
LZL2sAXFH6+6SB5LKVoRyxaFA9C6V6fqNVeT1yYuEeG+FvDDrY4JRtolemwc7Sn6nNBcnE5TfkIO
y2YkcwAPflYHIMjdXhQF4zT87UYhuEM3yLEFGlgg1C94HhPlh7GvTbCmZGXRt1U0r+seUIIHbgJW
9hB7pwd81Lyjz7vjdIS7MhU1T2/u9ySWmnnojBRxf2uMwCUL5Ytd3YSnwLYxDLyNaJjHWGuX7jUO
HBhDLha9HGdEosU8qp3EA4hkJoY5CBLZA94NMEBu5/UgV4u2u59C82zTbLMf+C6hbP7i+LAmkWlT
CXQvWGRxXqDgOg77tY221Rb1CuZyUvsBHoM/DyVCZYF7Tw2OTs+YST+1koknX9L2AJV8xjOOJB4K
5wuCxa3uJh3KUj03CLhu/pf+IEnlGf7t1mGPWoekIV9n3S0UGzbun+lUzONJJB0jPw+6NU6J1gBp
cXfbUd6/+93ELCxlRAZQ/czXwoqfS3Ld2dFWP3G/8hW9+S4I3l+HQHEtTUFvUBBSIArBNn7xuf44
tQe9Zf7Ro1biVy0ew2/bsKN+6pKEiF/iQRLhevP1Iog7TVJi6+6mzycihOHqPulQCUA0nV45XMDi
Gt3QIhupV7XV28YKaaUPaxBeKfnodXHS8cV2fu5bhVTMjINSm0eYs76p2+hFRX1PSmsNLTwkSuVW
wwxfvoSjSDVTPxJPMNgRxWYo82/k9lK3SQV3nNSAdDtM06yg89nq7wVwrBCXy7j17QhmZnWx/WQo
kqjAmyMGGcUB1rXKSfwE8ST+QLsKJ3fiBnZ6nLqL2q+0hP6Jn164HuIO+IbaHdkNCWA76Z87mVYb
z7Nna5Yx7pXztd2tx/GmEq3pTWBdq4O2d7vd8qLlofBmaVaRnM1AdvZiDNBvWVZgu7RM4pM1ItBK
zjStqrGw6iMIaN/XJuIzYhTMSyUm13Up9fIndbuHE+JoUkIpDARA4F7fogUqkDuJ18RShqLJWvlJ
aU4aPSxxRFHcRAoipDJWRTp8eSIjbk4LYkcQ59xQSK0s5VRWGVH5oEK7MHW9bqhE5bvptpXF5pDk
CFwcPd67DJgxmUlcEwYPiFyB2hUyKzBREj5SScKhifC4ivSx08+4qg4n2lVrEQ3L11GDhPLr4U8B
+6yjbr5UMflEdll1rNFaX4OAPPQRbpzOHFenuRLrx/QpApWNUmEubKVRjYiYfRyDNdfF3alJp9uI
YAvadOEfbLvP40pTNPY8dEPHZVjjCtO52iv9KKnRcz1P8rZ7d0o1MEDLb4wxlFKL11gOaPOmnluX
UKdE5qOLZ4WLYs3trMBT3BKjCKeyho4o0v9tp9d3xJRbQr+3e+B+lqhmPGSnKDRxCZO8+KpvnVh8
Nl61X8Sao5Dxh6moPgEe/LUFKolFku4h7Oz8i78D3LI5TfTpFd/J7k7p2s+/6Oy/AH3BPyTzBAYB
GTxJ8x64AOa9/1Sj6yDcx2vdLaDvCAHjNwF2oLMGDKM3Vr3/9TTtjK1q62diOSaeGHVLbfQOgZ5y
Yr8AWGREK2ry4Ysbofca8h89rmeF4tH12Ux6zRUrhJxisahRxnrUY/1/ZK6MYXlLrTKpyB0/jJMG
VYAoEC9xzxt10qlh/nXXSFcPbMBzl6EX+qAn4TS+gmhkHnF+0GTHtxd0guTaCr8JOD0e3BspqHOA
OOBCPWEcFP19YGHQjif3+y8eImP0oNM07/3yH9/Ly/67gDkY8xv/tzQ+0cIN2am7XhpP5S3EWEeV
2UPbl6YuCjURHbkkzk1bnddrtTDkvsTVY+ruCIzwxvv8gyh7ON8X/QfGWvo0TP7fX5+xRMUqTS6P
ItNS+dWrB4M0mgaajmxpKlwMyMNVc1QpalQhaRCDx5dHc8x/WhbPbRjX/gbVtsvL7f1pmg8LUyPm
Z+qpYoT4ICWF8mTjIB2d63ypUst1dn2WtnXuLGlFGsCt8B0sBe3TU0On071eRAcF+7U1iYro1v8G
brNLGkLeUmDCSOXKoAttVj9glV75XI+nMm4RXXGSXrPDqOLDCnqU8aCp3JSLqZbTgeURCMgiNYGN
K0Tn//en5EfasH7wfD4nIDjevytFq36HZjTjNUKyGGl0BkiMzv+Okbw0xVpYCF96Txpy5O3SWWEr
JC4tYPXg92YVcD+t5NuW5bSnuE15K7nRxDzku1ZbB9fK952gt1CYXxSAbTpoWmSb/04cQdSlEIeL
BLXe0MyCcFwTMMUYG8dirjtcyOX7pU+r1Hp8aa1wOrMWHh7cgBhfMjXY8dK7vBVaIyEEsGDBxput
pvYJUFLWGv9kBI/cJxp/c2Gc5pCvm3cET4j5Euz52AbU0A3g0/BEbBGerUW35smGUqb/+7sJXuDt
PdczBzUc/Ya+WSi9b4/60eR9z/Hc2CFUBADjfBEDFWbos2fiJpwsA729OEeNilBEgf7KwGR5+a8a
Gp0xWoAjd6eSWbhe0xt0xx0NBX1PzPt0BCP0Uhhq1YZjd7zRW8JscoNGAvMfF4DESDaB7RQM6sMe
5psGdTmqCL2BYFhXIUBAvBvK5LJ73tlf9AHDvgppbacwo1KA80CVzHOJ+UZ9jKXsU+ZftR6wSBsn
w55oCNRQbzOs8zdh7Gd7n97GFEaqhwqgCf/2pfggVX62bXMmLbXX6YjTtGCqhFVy6X9Z412Gp82E
nJiOoicJ31APvgUhYlnUCXB8NRJtsgAwj0XTbg4D8NXP8QrFJo8CwhNW9tdBQhbV4/VwsVI9tg8P
4jJB23ul7LKkU9NQ5UPsI+YjMWbsPaLs9pfSa0Qq+T3UxhE8CZsEWeMPLUxbUu7+XtPtVbxEMXru
5x0zk4UxhZK32+lO3qvHGkxWB9JM37ZwH76n9kmYOgXTFbgzLmEEJsCKt9cWtDw1/og2vgut5yif
fy5Na95/99vSgqXRT3e2Yc9KarXg5HWNpU6+fsKE8/z12fNDlso/MlmTLUl05EcLwCsQE0S1qwMH
mx2pMN2+VwJuJMbmZSB+rAKgXs64wJ5+K8rN/hei0MQXgENdhxkXZbHgZzZkzb8kAk1kqpFDdkyI
6xG5tKis8oyAyv4uEdh032rg1xgzCQQpCxzWO0eAj2AOnea4uN8zqcTK/TfqSvW0enCE37RF9yni
+Kc94cj4aLXMhu/u67hlf1UKalf6Z2WLPxKoVOyFwJSXZ0Rmpo+yBlYdy64WrBzStxDvxvd9yH+p
fHsupqJWCZKL55dvtWWXk8oFCmbMdGr6nffYDNIxgX03hMlRen36JQ1G1pj8EafbxKk7zTSFOewV
wCBsXLs48uaJZPQhGjCsXF0r2xil2qvBJVcVAm2FD7Y6o6ryjBEvU9fQlyqqsRhduY9fF1NU6SBA
QgYTXzZ1nKuBkf4XBSpQ59HZOEddWlYp6biT4wkC1a8XfFkV0u8MI9cfCXpB+VZ8gmTODhL46qt4
pnbaieqvQbQAseo0U+kU9uENQWWK/DPWpTIYNqiskQS/9NBlPlO7yZD+HkDfTM8qhVz5Te9M83jA
84WRQXrrqB3s+nNliW1oNH4WRfQMkCouqNRZUQlZ57val9Tej61GK/hLbDF6JCMRstjaujKyhSF3
4NgTfk+hTw1aWqkTt1+X348QCwoB7AM+3gjH4k9XwFRQUj1MuGFoAet4Z2sXhoaD5c5GpDCPPYSW
toQfKIqgM6Q1sG7138CGKUnpQk2tongChNQHgCy4AyQuWMR/VpzWIAmVDJoF4R2qk2mGvLZ6Zx6G
CI8LJo/0IDL5SkgY/XbCK2BGCvdImxfXrXM5QxbLL06eiHaTkiq/026VtpevyntRRwCEmvm74WbX
VR0tqDvWWyubc3aaNZ8WWqxaM9l+LZ9yzfc6vDqsyA/S9ZPlUhRlZNdhLeYwn/eetHAElaClexP6
5kJfMTLdZfeGSRE72KJ9uI0zmJ4GNWvcgCPf1dzPF+v4t9ydpS/rXzgrv+e6525op34MO3vAc9Ta
/UYcco/iSGeKy3Xl26cm33EESavhwsU2qED5wAiTOPM7BFjtgg4OE0whgGy2QvtoTHoCL5FYYHBu
Uh3/038Mb4VXy6S0EXSLGydlBEE+XfpW8eiPKq93LJwyjL1pzMRnPN6KX0X2AWELh7FAIWfclOGV
TXEiy2nBa7vzhORuH46t2US6/aLpoXAZ7EUyJqq9Y4l80pi9nUylGpXXphLogchKsIQ7BY8cXIDH
ACWfn7hx1sDJk+bCfl4jP1CQjmnRLrmylJ3JgSy7zVb1I3ijBDYnOrU/K9M89cpl1Shgy4EMCS2f
9md+Afy7z/fNFMFA8FPIrLpElPrUmO3a0zlPbjFiwVJyw35nPFqtzYrEqZ9VdcjeB16jsnZxpcuf
wtbwFoDkr6X8r/W9zGPfFe5L0eQGhOeatRdBu7eCKfeoJJcv1djbE7qSMrMklZAYAQRcm3aZQij8
CWdbu7K+XVrqEtmY+xYIOi3o7lS5NuT7IPmPRKAWkiORPbcFNfFp3L/2zWY1Jy/BxNEM4A5swtU7
xOikibvYdMRHCjVHhANOO14Z/9+hDm0hP2jqySv5GC0X293vg2EsX4tW126LpgX4YaE/mPkrXTls
de7gCmVGtZuNkYPmhzQd0V0D7eZ9vjDSBm51R1QBuQksPX+7tFeLc03Z0flsLC1x9ICu972ZGAnd
pn9AcGby/9OfYWVDd5iUZBim9ph3/JJPqLY0tRMkgErpnoBSCfTCsR0ij6HF+3Il3kQC0yGsPghD
VwNA25kYfLpwc+xXG2F3aVVx2bLgWoTUrnS79mnAxNjL+gg/eaSu+/8b+bnS3DY8SiQOxH8leziZ
TPiCxxuy98XG8Hj8VY7srgGqv9CyTNqRmg32s0zLiOAsOM/oJjjiG69M+lYcDmAPihKTzk12I7A7
4NQb9x0BorzuCtDIxdT+g7Yc9j3RqN9lZZAR3k9c7ntqka1O4cg9psSQLLC3LqwOJA5r3rbLj6xA
syd7hzTD3LtA9JA8+/5AHXdYchI9hjiwxWadEVthhRSIOhKAZi/Hye4Ew1qSZXfKD1dzVsritlTk
S3LF10axspHz2AQtbt6UrlLk8btCcq2Cim284ahIZb6ItXBLMKKGHvjE66EElhII4Fr1AG6KOtUV
WitZsyh31IYJfzA8Y9kYaT4fDs1ins3BuavtubgkOpMRQvJ8SJBki0bFYdUJsmgrMLNJUkfF+l+k
VuoQxA0edUV7rNLSPHs/mHQ2Irep08MLlyFfZ+YSymExE3R2csskMIXjg1ZnXieU8a8iJxjZj2TZ
YfDlfgWoj2rK9ThF46R1o5pSTJCgHGsc91EYVne3eU9mbkPyG/p67eg97JrF+uOvCOhW3i5aLNbD
mBjezgODBb0+WG5cSX6uYF+S9dmvTXQC1eAB8g0jkK5KHab5J63PNsTOw2mBVs8C9ZCp8Nkta4NF
bxdd5+0e2yGZvjBMmRtj58WEVMSc4BJ2Aywg3ro2WHt8J1tIWUuMXixV0t7kSowfFXuGgW4XvFzY
8KgCWcbHXk+62YVabX0leNbPN6+nrPJzYRvkzXMvljVN2S45zXE4mu983MaJNY6p+5NweuwfcPv7
IvEqdkIhCuFXmu3Y1glBOC2WMouV65Nqemp5fbAmAlQE165hP6II0S0aVav0X84nnXSlkyPYonXV
1HPvpj34XnDtjv0wd3OQxu9U18ezOGi3fq1E5zaVGY9cRz+vWsKji0o0rq82aGlO1sJlxMc0NAO1
3RND2AHGkqeo5rLyantfUnxpzCLp9MejD+hfJCTyoeHF7J7TlpljmGHr2t4tXac3vCPxqWLmqwDN
tz2mZehKUlOk/pmnybr5f+m8ON296hTStX2TFdtCcOrMUX5fw7LCTe9IbNUgmnmso/zbMAbaeidn
6ipKg9BGYKAiHiyMY6oDAFZtybGklVATPw5vP54strr9LiYQJUb6Kw/NV1dcSRlVtdTuF4uEYv9L
oQb40+FlZZfQg4ujnabZLMSK84iZfsV2jwQW4mLJlGu6/GvIWdA7mSMENxx3Ba+MzP1tPfb7otpN
RCuRVikwgqJD4V9Z18mzOBQMOFzSvt5ocLMu1cDktyG/bZYrQix4/H/F3W+LYRjXAk2MPPIbi7tZ
xuwSL39XVhUbBAWbjIc72j1YL/Nb2+V3CBeu1ZESi0xcwCer7c/Q1CYgnr7C/E04vDCYzXqfVKXC
UMCGZ5GNhNuRzSGvAFUS8QEgN89DGKcZQAxqiY62khCDCNFXhAprBjhZSStnEEXEGW2u6ojJUJwk
VKDjCzQlgrJxgfRTdkwIdECvsWmomtr3dKZuCvhm5wd6q0o1vlPLJwg3/0FXlZChHNS+JY1MtKHz
G1xWGDYm3VhiwC1Cl73QRvFYl8oSslp18puTBpfTJmxQqtVfQPZiVI/cOGTf2eQX+TpljZsa/WpZ
VnfNx353gPT0mysRBwQHDWtW3BSyKPZvJRPn37Ujmf83Q6nJXNLXgq3ItuRUxNzdKoACZCXsc2ub
7oaenjo1TBW50xBMGVE69AF9ohWIF4ZyqCYRvNme0guzU0XMAMFFlrOrxE9oWP1F+BgmdiSLPt3K
hhVxqR/9t6rNGzvY8BEvcKzHyjv7wlwN284exls6zImu+QTMgppTCJfj+0Nie/X55Y8jberIagkQ
lkZcBqOsEO5gjXe2k7znGhFxbX7la32gFWaSfjgY6YYODy9X5m5P/R2YKr2HKhCRXRuh1yxT6sV7
PJYrCe4AFCtgcFRG36fbnhCAt367Z2hOyEVxRIgueFaDywiUt9pCGUCc6h2sfx5kne34UBGRlGA4
2UENlV6gC17xTdqUjTy/w73WHcG6m5vXKGrQHzZR67zUp0suEHbGhgnHLxXvlI2oxt9qcSBTm0tc
v+HAdU52DHsiCcKhMVv490W5DNV3CblCyy21VPejbFY8j8PxQovgQlxPnbTCdOTzBsTkddSsL5ho
1IwjjyykbKP8Dxyjc0wBL2/alORC/vnWShxZM+UPi6e4x0AK6NWk4Z7GvP818EQuHBl/36dbwkgz
LNNudSEAkQTJuE0wq45r75TI1T2ccr56ssG9fq/RSUTkfbat3uXJyo7q2Kkmnz5+TnN4qF4UF2m6
IMflSa540ttMBx85w9c3hoFBSdcepQXBGVEWknHKW3Hw4ILDTyOOP2Yj7IcsMCth22+tJxhTwU4h
2eOk8oL91nlHMPnRdxYgKdQGy+0EwKe4JjcS3HHIMGFb8OE+yrmPBFOKk5sgc2QtWEqHnECrR2Qk
M7n1CghZjxrSkTM/1NcyA8fq7nlYAWhwJFYb7R8sGST0romD0nWmfXZiS+xBxZzHREPHgsTQH3la
zMir2tUu3YNAj/Dvb8BU5F2nlJQLji7VPaHEZU13q+qjPMiOxM2uL1bhta/Oq6M7CXHgOZepeH5/
v1ezB2UIM/u1LNKat9iKMzI5sZiYIzUUd/pLoVwFw8SIWhihp+Bq7bqyI+QHn+YOscGosszfuHQu
IRr51atDSPKlcnlqnVPS5bIU+hyCHVQ5cIeltmHaRtX85pu9lOgAFNMuwYGd7J+S2gWT0wBAQ6Ee
yejZjbdiqg7DNcR7sw7outEf8zQvnq6l55C969gm/y3mTmvpuJWsdV7wch0yYuDF8wuFbQziMvN6
qNaD2XEtPwkAbdd5x4GqTj/kvVypVctesc4wJ2sVYVi57g5YdTokG8EfU4E6P5QrgOcNCOZc16hi
d4+g73HtVsKfEIPC2Gu9u3YeHaL7HfmFR55/wDBH29ot0kn9OqmHizW8gFD35tHAZPEXRwh6LE42
P23ApnF8vWuO6qpt74HzwPgBkLNR/ruYAhUQU7riGojX6gyhsX/F8AtJn0ZisLAItathN7tlcicM
ldIlMTo1kKg/WpJ/n4Hi0SXI4VBLy54DpEo0rRhUlGWTc6bvcOKbEo2txSOIJUKc6V+wd7hQ/RBD
vicH2yW0grWY2TnLwtZc1mNTX4tCFoUXBLZeawgvhMIF+C3YS4SCFD5FmKmIY5gUrrCdJGGWe8zU
7+/12/O2sYrBlsfpMpSOJVPYznZZ9btVeepg7SyiE7ax6v/VMfVwJhGXhcHxYc+7g6IFRpEFHQDf
miyVHY+zhJ1YDQKqPjYLq63kz1pmfG47z2Jdy2GwR3gAEBKhNiWWbjIUBPefzTP7KDzPc6OKqc/N
Q4h9KeCXUAz5xH+JUTYQMg+xScLXpGuwTi8yH8L4W6j/1VVvUqrbqos1A9iej2aGKhvLXXRt2/PF
dYIONsir9OCRDL6XISEOqZ3a32SpLGR9K3utTjnqBmLjhYRuzJdknY06OTJbkdgO5ZybqxOGaMm8
rTkmM2kH2WoBMjQ5W3MwUxL/YBJd+HSd/sf8rYSVFbFuahdmxlrOTHhU8R4zBLT6NK7Vt0f99UgX
26HP2Cf7tz7CMy8eQUzL7aB1r03Dgx6S54ta0s7ldGOcyxHC7LKeKoGxVH1tovP75EWz2luNzVyl
qHs4OtK7B7Skuvx0jX1JQ3fGRPvpYSLkyYX25zZKUhdgPk15N6btFInOTlXLZJCNC+FlmhEApBvA
Y/zvK4NZ8zSdhZ/9ze+MhU0ZrDPsKBPJXUrrPhAk4KJLZxgYA6qdmjA4aqo0SCWPH3MzBJjZfOF2
VTh5vOpm3DBZadbhbyI80tHdAXywDx5BNy0/Fwjq3/sAHFoOr0oYNhYwfFMAHLdEWH58buJuUjVK
+FOPuszCRTc7LRdcfgX318FGFKUq/lSYkcVYbZRKa3EsdZoQb4agSV+GIwBT4ag581bxt9Ny4WBC
MNpcm9YMzv6cn58PR2qvL4CtEKBfuNVvUXMUXR4ZsJDF3Kp9wYhOpU732vE5QMdIR7g08/5j3+nH
d+n+FAX1FuhcoME6ESvXOsGq9REGx0txz6SDmn9YR3MQsgBMS0Cqy9tb1jzX6u0MdIHUGsktE/Fz
4tiCjG8N/2WC2SsW4p0T/m6sZ141MZeinj4PWHl5BwCHHnliWUByI5phkO0hY7evXkcWkYv2rYSB
yahxZ80ThG8dOpkTCpZTIsvf5sYX8ETaeQYN3MyRCt04n3WurFwE00Npf9TPqm0rh7VPGYX07vg3
rrBSDN2299q3yG694Fr1Mx8TKHkjakIjVoAA55nNgHxnAkLgRBVvyN8vCtAPy4nWvOPeNlU3r20w
uLFY8AREFYSAzBBFml2+rEoLKSf019476f5Nn/w0fiIt+AhdDA3Zr9ET9X+zdEg38f5E2LOH34vw
utZ9qH2Hf18Syibawlb7QlzHAa14oXoO2aZ346vAOmcZDkcR+Cupphc/tpKEVKAI+5MaTjlIqMKn
odrMvs/kKh6Bxox4HChzfj1BuCj7il+/W9hdfVhe012Dbpgb1wqCXVD8HuUuMlFOXgf/SNisFyxg
I2g/C9GgmuOeOdH5aUyIdx1cjDgxS7uK7044bvNuDhh5tZjUa4LfnC4uG8t2g613sD64Xn5YPVKO
lqfpG9ke7twPI12sraGzzxwxKzsc1Vt2iwtCWc1v7ABAesRqhlSqt+tmuwqzWMvbIFINvzq+t3Jw
iK7gEsUMkTvIX/FGF0oHAn8vIr8yD6z9wjxE8Ch5GA4jdfGkUdkSYWQid0heK1RsO0e008jJBRva
zkzgAcETdP2LgmMkCabzLWx886JtWqNeX/y7TvpOstCkN4RHQgGcIoqx0nB7FJFlfhogZY7GZjGl
NEhnxIh8ZV509zpcRxSQCvWNpVzVvHQ3dtXqXnU3Z/nl1Ogawgxvl7ZrQ9m2Fi0NagfiQ9TqFIUx
Fg2gWY/ehZm7Ff5l27sFIiKnwgqv2cRHglM5SdwQjdxexeSXNQXmNVArmDSPQ7RqBthPDbI2oobq
+zny0uJI4nSpHQy99vgwpZ/Q945a9DSAJzZxkxijM4JvbbeFXUaa6bGG/iEog08ubzi9VD/gEHGP
FTksuAt0c0lrPkh71eA/LiG6XDtGq39/2bEv1GS5b2OPDMpCcbjEbkVfXCcbD0r3ZoMEoI4/c6ye
awC1LITYITeZVXrdGJPQwRmbba4cPJUx3655EJosHtR7UTAgGw8CI1Zph1NzesTTw58C4uKvOxpJ
jVoNJyWqlrOyvFhmsnSwq9AYT5pB3Yttxckt27gNGwzIE/hViZ1V7jeheWk9bgSDJc+zQ6+Vxhob
BJmnDyrqdfQkIOFrFllv5ow/wlq1PI4RGwxaZ+Rd0/XfaYRhTmoaO3oZdLZULYeYeiqZmxJyOoiB
1aCbAPjHAa5kTRn82uHJICL1W6uAKuTefT5Q2gZwL/5TSDvjlqjBwWXYbE7I1PKbniIAv1BbuKTv
LlSooCchEhZujqodJ/NjsENxAgPiboJY/Uq2Kq0pNlG8/6wKJbtkeEFX/FFsSin81w7Y2RyuegtU
pSBhLm8Qmf7RbuZgGkeshG6Ex7VkCSngaq0ke0rN2Q488LEWQKlGDPgqmg/F/09XuRmek0t0YFk5
/hWE6g7nfQ37uoSLiE56p2WtLk7zuV6dFwT+LmIlf2fOjYLfKqTwpxCfS2VI4XN7BgvZmlmeyZfC
jNOtcPOC0WCEWJuGgMLFwVW0mleIWlhfxkx89lt6gQZ1ght19jH3idrPoNcEPPEno97zpbzgRvYt
h4aoczrOoI8vfZcO9mwJKXCtyqhx/gN8B1RyQ3WGY+/8mEaN+ZvtYpP9Orompp0gqSa0TNdLh9My
WVzgf7cOnU/YrceuiZGlzPo1Q6DrnTQrLh8/iywvXCdInYe9BYJPQ1GxZ3lXQWUBdnVhOB5e9hbz
jFxFbqzcUKCI0CUWiN8Zi/JXy/6XvrKRmmXmC5r5kwOkevQiBLTUjFY1E4EmC2GITE7SVsOMrOZ4
nHWhySVfYhtxFQxjpS4AQQ5pCzT8nq6wjwrDapgPbKbkCKXwwv4BMlv4tfOjpm5UBpnwz8M0rG8k
TpWAMCelXIJXIQlDF70VQVw1V2jluJstPtPN8CEYOlSQ/8tuvWbrqAEw0w2uk5+hY3Y3MmR+HW6B
/5P4XtIJVhhMM90HNOPuoSBGa0+ALPdfFHwC4ZxkXEa03uyx1Chd6lPS9czhPFPzThUdMlBVJ7so
v5F2DSsLDcPp2As7zRT+7MkcHwu0Af0Jwuo1M3ec53rDHIsbQ/mXz113klsZQIgUVPRxZVO8Rmrx
Hv6bR38qezdQwZkvKxi1yG31BGfZTGpyfrGpYsS0A3t/l7rYYSTysUdcKmk5uZ8TzAQWw7yxGfOO
yrXHY44L+37Pvca2FfmKf1Ddej5xQSxpn/EFVpbJK2BwfmZ2w2FKr3Wpw4oW1Yzpzgh1T7UPTRZg
t/CBFrU+9+xcn1LTseNmWT55KnGGVxT6aiFSGN0/PCILYyZ8EEVGcumq2Qud/4pdfCpooCEbKtT2
Dv42RRPKPUKQSucCWlQ+Rnt9jdOX9O7GLmkNDYNxmXiG98OgdYItGL95nluAq2YaTAlEld/Xw0eo
N0I8OPk7saG5DvvfghKAfKFQfc7Sv5ZyEx23BIOLY9Tbeeo3jsGeacgij89YWtI3v2/laD7gK4EW
wxEGkxoBMzLNIEMcWoOdGrYJrIixcZX88f17QqtJLSsak8zjDXiC0GnrQvX7PgrbGWIJ2fw512Hg
8kVyfn5gmz35epn+hxsUyX5UXGxSdgD6KFA4UamQ7bGHI6Z9UsW1wWRI/kfgoVIyBVmxlTx+sCz/
FxAEkgtlEYh4pdY2gfpH+dxQ3zpNsetINorqUb2oj5/DJFFAKYH7Fr8LqlBZfGqbHPY1iU9+afNW
u/vyxAE07iRqebQQUCYQZ8qLv5rdcS5fkpZ8xIdQ5pfnV1BpE3ybeEVkn9ef9NPWKk8PWPjYnmcN
SbvlJcaDqlGKEq1e9jbXU3akJStQmFQEPsgW8lyHBy529X6X7xOEz7wz1cr8YRIX9QgfTCuZHP6V
p+tKjQovgnpiPb8j4pwyM+uCQWEWeHnhvMigIiL093xD0NKcsIWxSx8ihvb7VU0QqzHOIJbpd3VH
56KGgx6tdSDc8PXHldj9t0HLUAzGQ+lHxxDYm1TEEDKY5PYFUFnvJq4B57uPqFQ/RC4mv1vl5CVD
hNgA4kEUcDX0rgSE8Sje/QeYZKH/hmoccbp61zLRAcrJbWy8YvxSeZ4PF6vaVGoS0IQgln1O0gVi
8Dp0T25CybF3jkNAkBOCaCoPgTli73WhthxS1LVwhuZd2mytlsHzzmnxnp/Pw7leFDmThfWVYcZo
DYnUIASZ1ZvsSstV+rjRDGR/MPs8BxgI3TTeIlBHN3/cLbd9pxW+kwLi9SPyopJ8l+NArd51nnu8
+jMJSWuO7Iq2RpHgbm92z1AKH/d0m4ls5k6kPxSRxQFSYYLlz8yX0e9fOkGadKFCnPTM9i3YWNd3
Xrc3lzCCAHA/5ttIm4bpDZbjNu3xquoLIVXtSzgKVbJHeo/kMxcda5E4D8S255QeQki3FeRagWQR
GmUnVayo87OuydACrWrby/prvueOSXyDK1SVXmd+lWOgTWt8GJhrkjMwD69zlG/YVyrTCqiqrQgE
GnLCb22ssimhneLsFWCzG1r/4Ylv7fAYsJW+W/9w4BiinBeASBlfQ2VrRbxT7kdpCaqv6gKqyu49
iEUTBZXTxBOOaTwCZzFbava23dkqti5G2IErXwZepvQ6Q2Jn75//Os3psRo+BGG5XoG1bhii0+dM
CmMYP9MzkSTiRDIVYOZT0QJln7yH7buOIpP3pSzrKws6y2KVWY8QVVUSpmJ40Ae+IGL3Bt6N0gKk
uXiXxq+7WKblMwnAYDXHqRmxYpwUon6MQbP9x3CxA9ferU9/D9Vs/McOV4N4GZmiTGDDXAYFFJq/
3ZF7YsWJ25gjBUY+eaZBfwgyLiRp3Kc/4W0Xoc/tjsOEUQzIaQ2sb8Xy7eJpnAOWbc6GTvVTAvjG
gHdrjKfpU7SLpcwmrUwHs+ICZNtIhuyCiGopNO0Dn/rh9QVR87KMhynunarruKpV0XJzfKLPB2TR
ywkofIf1omP9lxEnkkISO3F3rKKcxtqp72VmZmvehwxZZjeCqxkh3gkDQMaKelLL8Cd2H9HCZCm2
pnCdef8la7y7hmiUD883yvw/gxL4N+8Ft4BugH/hprK6oTctDTiBReS42X7s/oYv6gu0QJdKPa64
4lvz9vNOUOitbJMMCMGodw9v70PVSLA6GHdV3b7PtiLMlJ8yv27xWP7BpMYpq49Q/CvlIMugOeqv
sXu/hsHeZdTpKH2bl2uRq+fmtFPZY3DJD6u5WROA7yrwqbRBVfFA/YNrNM3TM3j+6N1+yiUY3j55
32mf3YLwxI6l8CQueL7XmLmAVk1GuTXE0H3eupem7pKbypC7r3qaWtS9uyq7yDybwLtoeJunHo0d
Ns8dAvHq6mGbHNff/R9mrSBTgVZkd+NNEBQ42VCwcldni2/4tZpejx1j9mEeX04c8I4qQ87l3ev+
rFej9QGiQ4vv3PbmgPxTBym7Y4t2V6hqkcZtHAPFwvsvTA8Q5UvRJjHX/RAZM6GiRO6jcXRlQKq0
BSFhXmViOVCOTu+cWLo25X0EnxlSOxVnd5wHT4pHzDtUlaV6jumS4fnqQusxehAbrT/eyYmKF27U
qMyG4pqR+zPlJkFp/TfHwKujJ+0TdJtDCfID+x5+b3kGRFWitDYsnJ4RfWv/GR4Quujr/XWCZaLD
iNVb7G18drh+YxmnCtIOjYWkwEiWGfO8SlFZV1NKRnjZ/QCxcdOJZ0REbIvnBt7YOJwxEeXMusn0
WAXJmTOKH5i4H95j+tcJb6ri3bT49lUXUYzvoljH47W4DjycR7y5Zj1Tss1cF6Lllp6bjCnR3eh3
Bt+TsJht8xB9CGRsgh3jO9D0LdRjEm8DPgbzG+Oi7hMPQsivNiuDyco2GEz9eGqTBazD4QvX3H16
QhgDYOsuvQZfgOQAzqwRXwABv5Ug3HVCC2eogDiQHCoIJF01Ey0D8V4tLLeTivI4wmXJjrEZOBMe
RWHhf5axlk4IF88w+bqLEPmlhoXc54WRUa+YzeDhslsWlDZOnQLG2rFono6tSdw8FrAAGc+RhAuF
mlYZgPGbBzo71TSgG/VYMfrvNML4LPrZjksdk86jPDm8rjGOxbZFVSxePWejpdtI1pDI1seFDz7g
Zz8cmkOgbvfMDWY1q2YGbanwtbE7GFkm/b+ToO55FB+/Vjjy1RszYpr3J9tEeLKmd3wrP85eFlIG
24L6716ZqCFmEzmFPbP+vYJ9AYiXpWOxCUVCgbatL7RqCxbWqJVYHDW7RpffPektGGLmd9qSS5mv
qGKhKjA1UsEh1PAt1XQ1KSu86HJDUBGsu8sIAWyzCA3RYsVFDdvKQOIsbwInIVBctgpIE8YoJJPY
J+LEn0crm9Kqt/8B50WRV50gwm9YFjfxuAf1tiwEm6hRQebFilgaRuYg4diN4/ZM0T9sC2ciJ4BT
6b7R2zshs3QAn48dq7Yi59AWTI6K+BRHIjC/OeMjJ84c17w5gzdUQuxEEe81yolCOBi27ECcmXbW
7QKCp1m+fOjyA5io+htzYhQ+QjHPo9kBaVGU1Z3psx1g3JXsjKqEgldGGgBu0mxosqzOQTSgnsyv
N+mmG6auUnPTYJyXFluOH5HFjSz1JurgmlA3J6LxAAHxH9C828f8W8ha8l6isWyMusFmUuE+rhdL
jLq5x47xBb/FHoB20c5l5T2rItjNq51SkH1uqopqsU22LMCJVD/45AaAt4964fdAWQTklVykY1QE
ll/oV6z9/1NaTjQTwHLv5/zuOu7/QyDN0Jj2YZAb2qbIxV/qs4sC9qvfOsKlPToRX2btyIRdGFS+
otoc2CTgHa/7ZDGa+vZEbZWVoq21FRXQ9zr8d+qNdgHVe3Z7S1PEAynEU7INxoF4o7lAN9noSiLN
P7mEjs9d09wdocV4z0vkGTj8GbrsLl0WDPfNL+SjRDr8ZY0tam0m80luKc/VvyoXRrwHJogBdj3h
3YucIaJdPVTP3AIsatV0ozXcOIuXMxeuQIorlir0MyECEg7MO9P0M0bdVlPdy2kRhgypsuMw7Llh
AnPtl9hYWV0bIhIpNq++2WDqdahWVQaiMBekKBUtDY2GmTByGbpUGmC8XU5AGSMe1bbhWzV1x5YF
O+1rsR+U4/mIPgZGrjPZtTWip7MYMsgzZ9MYGt6g1bYqOPXvbF1vlAxaAOZ5l6xze1Ev2cij/UFl
mZ8EYobo7+5IGAc98qfHI2LP7Bh6nbeKvXFyf3tpIEQwN9VA1jAZtsWLYA6mxlrhM9xIZ3XkGBC8
DMuxoMu1/kMsTZoy7Td+gnhC9Z+YM/AvQ4FTYw/dPrJqYJDEswmdulb1Phfabi/l2h0FRMkfAAzW
75ssAaVXxOefejEP18u+xjFrkTroInRBeqxpUW9YVX4Fmcq5zH4xM03fsf0UMymzKbf5xnZho/Y2
o94RMXJu8QNEMt1TS1DXqSS7Pgnl9RguOCCRqeXp2px8B8E0D7rTeUCDdw2BjmTFZ/3gGMBvVedd
9AFb1DdvFq7Boc16bF3aglNBBZUg4YeKGg+YNACFQpq0mYvG1+O+/+4KxWiH5V8qKXQz4VV2WDQV
oNlO6pgxxSukslDjb56Kszem64dI3jrVRFFKzkkFDbUbJnmlKGPrYpM8GegwTg+t5AT1/n+UovD+
fwR//fu96rDlLzzzH3We5jGi/HDy/qIix1n/VgcA4/bEU7CNWSi36/RRVdJAnBMcg/Rvhww4Rv4D
o2GKXwWl4DG/LxTIk19l3y6ssIdqdT0r1GQWHimcksFtGddcP13rROwgEQekTtahyXSWoToRtJ2X
CrbXpxKXbTVNmjTz9ymDb4HBrCii1L0dnREuGIwrQIvMg968O3VJDQzNXC9vR3j4dmhwLFfnBwb8
UEvUcxgQwrY1rxAZaGWmumo6HD8TbucN7KxYTkKk3xGUXT6yq3c9UE9mkm/1Bm25BThdSNwUDBrZ
ago/kKqWbD19JG55mjsO3cic7c7wLWu4XWS8vdDEuZ4ee6zprE+VNOdYLgWqL97Ps89yyrOc3yp2
h2sMwIpIFuNnm911a6/IhcLHY9DyxKp47N9EMlHti7n/xwbSfnf8Q2qaqPTtrZuqrzxHqaSTZBjm
4RgJSjIVB32N50TKz+O0YtaoBulYnfGrLsEeKURQsb5J068w50hjQQ7kYRZSiUgqK+ikeYMuEGIa
3fTNK3iG6xrSgDYl6Exr/y1i7CGmOQmKa7S5jclEMaqu9IsvF/3CL8Xw0/Yh604q6NyhjaWCIvmY
59W4ny4hiuqeh00EkpjdBekCj85JCRnkIIWoBV9ups/zf1yEVvSXO4+NEpEXZhwzyNBIJBK9zot6
C2QrGAXgcJ9mAcRbeAh7ITdHAbaaD+wH5R/ZeDmE7BnvaI72FZITsf/wV6lpeQ77uCZFuxqyDMeL
lKHmp5qq4K03dSpg4tyJjVNaOPD38MtpqOkL/NL2MQviaeqWWhNtAv0hniuWT2Cb2EvSUqX334qO
2Flk5iMUN/R9Q92zVR1ZqU/21wlezPZQPclvD2WCFXJuX9QER9bsFVuBoPivXil0O4KsgrFt1rCG
TWyGTm0FyAAGJki37wmPxueQ5lrmAZwF7niOOwu4gGmDpJHtTxN3qA03/R1raZAgAJI+tBOozGa2
YIUZ+pxBH8LUsYC1rjGehpbc0AjbFsLHbZmCaxVsCRLwhJQTQpc5CAbJC0Qm8J6Iyy+6sWw6PM1N
f15X3KImZUQ4y1alW6AqhlgMMqnb5CF4Q2hzHSeepWGlAe/d6ESHH7+3zPdpormaDJAvrdXzhSAh
7I6cD7DAvocDhV06oZ9E22zaHMK5CEdA4SginbRdcSe4S+53hTL7E34skLYIVREiYWydIaGzmbIt
u3p6NJAzArPNqy8u/hlxT3d+8lyjrJn8b679JocbWRFqDonAnv+OTvA1MkLN/6MhfRcdOCdHs9F3
WAIIK99MHuPw/2A4gGzEj3yP8jejMzvIoEF12nRvB72Ni/Ee9yhhcneLBF5LPosyCCprcRSuSH0p
K/RjSq0/0sKfymc8DKkpuRKuJ4pj/lyAQZeq9bGTWsJJ19Rrev3VICNSoZVIeawpJTDHwuBaxAP/
GvpqNfQEyTUM5DlRG8up5ohMhvGooF7wrrN8JRuSOvbC7arD/VqBevmVCryMliDfX7MTn2Av9lxE
rJfxXfBuxgxe6IWIx+zE80aEDS50dbbTvTbvi6qdnjBAHSfrNaG+7KhETQLBtn3pN0Cn8oYo+jsH
MQ1R6Fdwg5+DMUpxa5SuXB3GDjWqP+av5RPozKA8z545Vihu69YwZKpSduOi65kSxcwUCVbrIQ+K
6aTS+ap+rjoXQP8lVVzw1AdoDPalaM07pvUvfvAWGioqHxnyMKE3BSiN75NawdY3YrVxbS31vdXg
dMPFI1CH/iBe3XSAseNXSQLqVWf71SvzrRVJdrZapt3rUGOiDlXOxRHV/qXEgIo+oXtI9xRVQlJo
kkLRsnmugPq1HaPT3Qu/Xeub5mmjBrt1UNe3LieDmP0z7jzvHrV7Nyne2MFTeOaJ5WaZ2D2x5P6f
3iMsMjZSSipi06RCAUbBBekfqI/I/kbZyMxJCTyWRJF//3QKGcW16vqpFdAu2RsMFgLq8d5pE5T4
k5FxfXnyT+KGIO/I7RvddoBLihkAkJcwBNzGr/wplUhrvfcxqPPC/9gbj64JccBGU+J/0HmNWhup
m+4nZoG+c0qsWHv6WZxwZHki6L6xP+Y2u6bjLIr4VAElETCRkgIhq2009T0nl6Aau3s2MdgmOWCM
miEpXEUTnD+3KQSsqyWDAqOR89M6S1FwRnLwmKpV3v6nM4PrTjce2o6MO294rVM/YOtcfgiWRto4
aHsyPK5dJpzrGMn3WF/cxFsSIT4LtD3GrIaQtY+f1xDSuu5toNZM6hUXSSA8jed2BS8B6UsZ59Lg
zQmUEmR35M14/EdgsOeNeCU1KVOB4QmmCuFZSe5YtI+zIfmn4zmCSxjlWuUeuoxBBZcuE1+l9Of9
vq2wwaK0LfNTcFRkU9wXVZ5yfQ4z/oaGKWJ3ba7JLTkddNi7XBfE7T0wVlob7VS0+tFp24ZOvs1M
d3pbIbH8k1p4/NbRcdnhnGYJt1kAMRAQ6QRJ82oEg+4gkwYtbF7OHFGwcxPFCvZ/R2RLLCdNcacf
QnXA3RTn6oai/VlWPQ1r+/3bvvSpY29MHSzR8Tbjospvvqxyyp2ZKWXCyqoleXnMCGilknDTZBOQ
tIbziPZ8lHeg/ukkLtR3SywtbCuAjzZWU125+7sihVix89e0Bfhv865YbgyKFLcpPlUxlUf4KMre
gfYu8gkaYzC3iF1R7LOePFjJZvv3/MSqJ5V0vm7MXdevfDpjjIv2ZA2kRDHOJxqXA+BeSGyNKnq5
b8lKfJrgT5XXMnu5Dcjs+UkQtguX1u8dudnKVcnCd3fY4U7l5IxSBCInSQ+VZKWq/hNBvHiFhX3E
rPB4B605CFywNfulqrki1MPY5JrIrT/Iq+IrSAmVQ/4TAdrc+rCYvxXStTEMm9AhACP4DSFoLc+8
WsEasQvM4XNjtyvds8Ulz/E9+okFnQItTYzR0ikPgpYwUojEeNjZHbq0AX0AtKtvbJcL2CawbruG
zrUYE7IYoeQaK0KBnjzZwK9aRES4dxylSeCFGOBX1nECkN1HuM480X7vWrXnwnmp3gIChy0LAyAX
8jhSEU4SbB6gff5hJlMfoUBEoBRk6iRCG8DvPPqp8vKvZJVv0z7cIymXsTbS3mfhCJx3703pqv6L
wRW2eUG0V88fOo7ORjBFuBunVxvFWGQOn/jLSmXBIgdcGd2wP0XzANPSGXOEn9a4nA10bskh2HAw
f/KsDi+Ezf7G5ESL1YYEW1mWM6C7AeO1xGDjkp8Oc00A99K6MzygvwatngEEnDtiTOw3pcUhqkU5
EsiYHGXA6Lva8i6y3ETrGqbuNP6PTq8B/VQrxwGgn1q7SmXeRxFKNhbOzspJVy357wQTPunUW8vB
dsGrd5cIH6HAclhQe2YhikB8bisTnwq9JKqEM66LjsrR5nvUJW+zxwpMYIplQ49DHMpUPgV3eX7q
p7S6DoKFEoQDeSNLpmRzBVuHT3Wl4NrAsHg77IsN0BBjKrhX4Morhgl5L+CpgkApVLu0Y71tjwh5
xYEY7U9gTnfd0nQHGvL7Sn/tY2UNH2EkY+ljtfrhYpl3SH3kMyfo8wHjcdFWb2Z0ZC0aKw8/GjxQ
AShugujNOjkvEyhUPnPtkp16Imkm6zm5XHwCSveFa7/esL0z5ZIf2uVgjc8oxrGLkHj6qfsDrSx8
CcBYA+RB8LUFwa96b2XOzXzSZXRUHk8MLK7iy+sARc9uWDKNIHf/HT4z+AzLjSQpNR9VDqx/gVGh
rgfosro4xd8fxIv4SIsrmxMAfnMP0W+eRL+fvin/+GNCxbR0QruLxL+ypSRVDpYDDmGReOUXj4xr
RnXFXRSbhIRmttzX46nK+1h7Y8H67t4MSTCqImAX34YUG2AaUx6N6XwXr5giwf61O/ROynZG0zrd
i8LuHK9nuY6DfxOKSMwNK1Rhd0qjviipl3EJDNXV3fPjAfFO1kCpqWCUc3tg9bD8VUtPHOa3Rg0/
InqgCIoiSJINhNCeqG/j5J/zexe8J6opckG1UAnO/TmbX82st4oqCpk6kfeSMku3EXBbk8L3tKyG
cEJfDDX5eCffBFIcMfdF19p7DtOU4A3Nm2UK1f/WJ13q9coQsECMHuBYUikG7xo4eAnp2NtWCZmL
tJBJrL2pMCj0UdoHuqt1f2813+TwcxFGimV0qZrM1w9y1VV4CevcDgwMGwzGVGANxbrjoGv9W2Qq
OtsGE83SEnN+1oRjUL/7h4vQFuznRaDWBvVnyxFTaMNXxfYcqOTDAQMx3ZoMQd+KoFp9YQuCxL42
GQkMTQAj2m8ON75Ox5Er6v9X1h8IH7KyRv5tNWX4idS+dWMPIvLE2lWeFP03ohmNtvA3bkqw2ZM2
0UwOJN2JaEMi3+tdPFVlooqHIQgoJB3YJ6wUBHUMFYu7K7HLijiAO1fws88Wtd09IVtd1BGFQP+3
TtZrH9bfZ0cI3ngeTmPmFgaBkRRKPgBNOvhJgQ6XV7SyC9tQakfmD7jcC5ThOWrLKF5yu8uxtbGS
cSyM5qCiznYTplxoDBvlcZ2xkTXi+QNGcA+vDNSmNXFa6imQLcaO5jR+jVMrKrupbtgS4M9A7iDN
uwn+xhh2NwLOzEoBN3m0hqPQai6l3/PsinRqJhMR+XyCbTn3czUUxWl5dAl5nIEmOPKPe28abmr9
acjJMEsWnXEbakCl1vxzSHsaV1BUzYzTiiOHAVLCM5irCHei31aAjdaYIXyevB23ktDooaCRjBUp
Da0n+/jBX3Owv7uAxYcmZI9ZLYFf8Ce4wrDynhoTAkpf4yh2K0/XeM5FiR5N7W78OR1E2La/5BKn
NiQL/iXU2ZEOJrwF7nbrO+1i/BlsvEA7SzfKjKmEILk5FiZ06/Ba8KZZ4K0fI/ttqHFAFysoskr4
EUhOCPVdu/l8/Evug3/YvUv4q72J9fYcRVrGDLVgDkUdLMzZbWu0mI9f/KWlPCE8iv9sRxmc3RXQ
Jay+/tIN0xbM67K35ymcCBJvMjlr2Hwir5ZX5r5/onNMRFYVQUiy/+5rn7dFZhR0HrP9CwDzwrGz
9+0GS9HZS13G6WmLdI63w+F8KXv6p/qcdyo8iVZLAJQuHWwoVEQ/rsdhKWxR6CQxp+iOFOCMXn1h
oUoWJnann20b5MxZA6oZ5aZe2+nikxP3YtcHut/6VFLp0b4b/rDeJKje7pppJKFdDEXtP9+aJXAg
0B/c4wjw/d/1xI7eFhqQ5TG7kFydhvmlOVb799oVALWkuo/tIT4+XARJIWNQqLAfO0YYDwshMzIj
UQUvOSCvmxD1Wm2Z2SFmPRR5qMAGtzxpDlubpuuiwVYfpoT7IkkeiuxAztQPbwzU4GmUyxvWJYwF
tcV8YaznPCExDqehwQeneYxbXfenpoMbtopMAnwzmyetD2pTz9sfDlDfj4o832fGFa0QE6o6FQVQ
1PL/wgHylu3YoRnadyrL+ouHDfFDlDQY3fmyagWGENYcJv/eLy+7fS3wd1q3DmOq3KzlUzxzC1TY
IML3bQstTaqdjYnMaKNyVr7epxdNlpbXGLKmxX7LYD5cYeNEFw+qSXZ0eCX38ydULSscb8Llde3r
1dkTHyygOr58JZWVOeIfmekV+icNb8L2bhXRjMONi7ppW1IB/aXDJJRQ7Gvjaa8ViXIuLf1ttKcP
9YVpdPeUDK01egL/30ulzgfTYyGHzLDTjgjRBw8SG6RakpgDAUJhKNX5nrtfvR8ZfWxsAMfenLkK
uIU4yGEph0apcfWqOvkgCV7/LW2IgwLLzmxXE8jAN1wbv8F4T9Qa+5JDRjjItF/prji8MDZFB0+W
1K2jnRcq2N30Dt8OglQSBPK5AAWCe5UZxC0NwLXnVSrYMIrz6+WWKNGAYZ2c1JMAzDdsqRd1x18i
onw3a0hYlTbCrCTWzCAKMd2T/XnO/L8ORYg6UkgBH8wMNH8lBOYuYg+hXTVYbHtHDzaRrTyyE/Wp
BUfNamkvvXdNfJEOL6jcMRRrRL7Ie10VPrx/AO+a1/5WpNPOZrg3/fpY14FMDU86Lf0xks5p0sn9
Z2vf+fuhC3F0dfyDOzoF43Xhg8hkNdVq7oVv10xLvlqmwn2LsQoMBjEpmFUw/KbQFoYsRhLVa/mH
/sfeRedVDrBVYmQSTsU6hWvO06VZrwxcnatxgfv0WHwu4AH/71y6hNQWm+6Mf8JM6o0/MvRCDTRT
GubDwtczSWeY9xjD0DGAL2UafTVCRgk1OjPkWUnBokExeDO1BzEJIROIx+4kGB3nlKBLsPfrlXV0
FwIuWjJImfphliHGDRmX/szd23FE3palS/lwWRzCLyuDXU6UyOPO8JBmda9rc8OhEQyntX4O9AM2
kehZF9PpfMPG0ItVgNuuP2xRtMEzCqyTnK9hgrpG7UjDLiqer0G5HmN+6E3sg6rzO9s7jFCxoQaR
kMxyY9ylZSLLec3ij14ztaaVfghpc5Q48riNWjSFQsxGWxOfF3nx85kXyrSY5YOttBKCjVkZjwyc
+EFphwOdR1bfvZWe3pw+bvcNLtDeZ1Fp6z/0vRvpS8fAnSw0Qy/+bRbUpfHYz9nh2rFI8XlDaq2K
v9r/ioatLz1JerEc547XZrwrqNVhVLDTL6Rzg2Dc27t16wX9rYpK8choUeJPEeY7J0J2oiN62nIi
0+/0e6j5nlo2NWvrJwnNTET8OPyE8I4e2q51YREuaGgYNPQjvBrzAawpRoOGkWpqdN2rBFrEXRAf
9uN8m6y4BNDOlTYu08z4BS6sFKpTCUq4KHDB0Gta5dX4ElV06fUkZrgjjCZN81CRtcNrYh1nhjer
jHpd05zQ+2DSnPmdDCe5snksnAIkqBt9QZpTJ6eX5F7R2QotHDfWq3ZbicEA4a6clz/leiWCAXUc
/OuLqqtNCgOimdyKbhdJat6EeYuFg+HPEmL/lzMy1qrenT9/dWSbH7zr6JglVZ+kPjL6yNvFAg5T
RODd7lnVkwkfyq8tUOk6ES4i9nh6QA37uaAdPxAM1MLr++YcEDCgYPwobgzRhWkdw98n6Wo9u/kw
DHp467d+5W8wSDMd+liyPZGaowuSWCIm+SXG3ybze2RPWCJpkN6nYHMTy+ryaQ422b9xBoo4Q4mk
We3x8MnQ45R+7x6HgXi3Zuckk7C5tgWNdWSaIpKjdFCStJZwe8wrAuinEmzxRuIQFQ2uBJfpRC3h
SsRgeFmbNIXEwCvP7zmBAyzmbcxz+H9TUZOsJM2+307YwiLREaqB+atooDi7SdmctQ2EjdRDGCUl
GTBX0qJnd4m89qwb2g6bWZJfq6ny7L9HypzsPRZcABUwTvWVTp1VLJKvXLauQATKljFoECt9hpKQ
zshxFL5+ZStPil3113xFQRDqovkkT0cT0VJX3lJEbx4eOF9LlQGLqNbHFoiOSYxhqfOZkXEkztgC
bNFZ/qPtOSI5h3kz/GNP3ibXW1OBKnV87PAIsGNWbUyxvBVJoK4iarXwYUL3x0dqZv+gBtJ4nOaP
pSgwf0Y7eEPF/JtkL0XbJzPey15STrfIIVYgK2zwNejpaJEAodb3eyqXJ3wrziQBoW1Sy1Ob0Faj
RKIsuhkplW0gBuvDl/eLHDtzt1OxeqjH5fMAG1uozSysoPjFCoqAeccg6ATSot7OBd6dULI5bNMV
Mn1Kj8/pQ9zmidppPXChcibZGplcIAMtkt1dZxD109KWC60DVIHsgHZVAzIxAUVw7YMhVhkgBN/L
zCr3B4knYD/Mb1NFhC4g9POwZviWz6AGnMMytwqLCUw4vA/t4exn96b2iuqPGBzuXyCrcpU/+cTp
BX8BcBUvfH45hgPUPyWWrSullWf/2VglMgETf6Z71+V3Yx9RBVTe2MnbUlZXHZcHCnTaJF1JUaAH
fyeJtSqX0sTddAHBjF2LAVANEcdeNSvEp2QfEaaZRd+Bi67dw8Vtce/0K2SlEpZBgFpAZutMVHAn
nytyFxKinPXPz/B1X9rmSfkjRoQK2iw2hgBW571Gp9LKnN/55DEfarxuXBhtGe1sVFifk7oKt3cM
mZ9cQDSr4oX+FoIBQK8rJAphpiR3rvYujLyOn5idGzd8rOgnj+Vn96cgu6SrH2L2S9n/YTaf8kl5
YPPvd65oE9npaJ6Sbm2VL96HM2Cx+rC7ABVWTv6MB/uYKYTO2nufpw2fnR4ScRbRWpatCRfKP0I5
4mBmpfbIEVN1vbvOUj6hL1/zOulBsH4cXfnqKhOi2k1u6kqw+JPWwbVF2zUHhCtHlEti4mjBJcq8
zNR6fyP3agQBfQ1dKcg5m8GKk2cQm2K8MqxzAETrd2jww+WERe93H56roQfNEegr53FYaCs7v+zi
X34uuKFL5K3Ymjd81zSScTyJbLprNj7W4eI+l54+fK/dqYnfYylXVKBPCLXQlSJNaZ0P1qaWfqGa
dFkz5iIC1m+TjI7+PaKN2WyOKaIYeQr7CFfIVmcX6H6aMLspW45SRC+LIWjZ8QdFzSLTLPvjViN8
3bUn01TPpIOM3JKCWap8hHj2LRc5xVeD6UEx1DpIgEQ52oahqN91Wzy5yzDBGz2ls9t9LdwGedrw
ewu878UNc99Qs/BWII2DL0LXUgPsOwVnPTRb3ErQIeR4fnCjAzNvzd5Awz8vUBm5vrP8M05apsGH
5E+34wB2h85t6zAFCBlFurdLvlMiNgYFZYAG8O0imG+dfEtGODPrndoXqmqSCZiLNkDRPBD2sIQz
w/y1n3xvQZ/4+eAg/RZElb/+nlbZ3ug0/Bx/nZQykyknLb5/mQoiBw4XVZhxoMp5fPFIY3C94ZT7
v2PgR55yaLJfeSRkT3QkH0cXQisiAi/mKlceaT4x0AoVjYKP6MkoWpYAjmQbxO1/Z/htbi/d4rE+
R/w0q0hInW606RZfu/CWixcpaS4Q/oRfd8ZcNhRBJo3yS3WXHTzP1rSoK7AAgQjqwsJliHy2iOTZ
swb2M0HspSMe+yJOVdJNyaYF7H0UsftHNu+CviFlDISPTn08ZZSqSwlHoz+tLlF36yXBFJ06NAoM
Qkf+yOreJKFGaarqbsJ1cRrJ0Yjm4WcgJ6BRVBOgKISXjVQrjr5PdEViwWr5ThEZz2qftG5KZEGU
dYbemkr2aH5vdkPs5rB7YPZhTE/qKLkddvaa6MySb18XfYOGM2qpfpcu0Jqki9OwStehVTO0brJN
k3t6o34c05tYzTuTsgh3UrE1FybrWKcZtbLoWEe/dDWdrWwNSmbXqbC+rC7BTtD48c2EmhqBnafc
XkoESG803D0vZnZNgmdYsfEAcLxTtH2jHenAjgBmqFrIr0WxgxDlfU7EUVPhh6HuIl1XBr2Iu7Mb
3g/DjdGvbQcdLgdBJKMtwnwexDWZDBS5SZF8QBfi7gGa9Zu+xopnMV9UyBg2zxgFG7mi/zYgroGx
3AcG6X4hLtpuLWGghYW0rQmWj30ZAG/JwKjleaeR5ciLRqc0+UhczAJwCPiI7+keVzZQ+O+e7IcR
HousbMuPnCfqtkuIyyEP83gUyhX3QNHGxRh4KdLyHIANuIMlYQXm9ooqxdxe7m+XPbkA0tP+PFQz
XdtSXxXKRNgbQkFBYZl6nJZl11i7KvAVfGJFwpRagZZ7/i5F11Q7Uqdwk6vHngtjxM+8oOVgT9lk
dn5c+aMJ/T6MylQVOi5ztmuBeIyxK5NgLoedlTqxeFriseevNnEBtmgTYUaBQXQ5dN9zWvpG0R4G
R1pAlHae7hKt9Pszj9wIBvelbdBLTBzX1GRnxzRo0ArbzS21J27UMiPZ2GcYVn94evJJ7L55x7qJ
WK8gbgI0wGTueDjtZDfEQdty34n4YCyZ9AEKlnh/hiCb6zytQlAI7q9+/2LljeEwcaNSarinsXwq
JMxhNOXhUHBMBxkSCX160N+3ppWmmcBdeaAXnANMJk5+eib9m6KYEeA2l++Ribb0rqFxmZDiUDPx
AlgK6MbzOfJPTn/qJF1fv7+RoJREl/dQp1U/z/C7KxL870yrzZ6z5kjyA+AKPwnsqN7ufdz7PZ8s
sa+R2b5/nyeu9RmnKaJNq7bQsm8FGINom4Ml6eklOW6Ao4+RTXjbtCKA/qlxnKodTXTa9QWkEYpZ
0fFltUsEP531wFA/IThurkxOM4xkh7pMG5huch8JTfiXBfzP6b2Baf1/UH2ip1dWuknJsclVfUhw
DXqufqM1idIvzPjbeloaqW9CcOsaztRaxDPlUmvdlo6dmrbXb6wFaR34ELN5e0F4fuarT4plmuUz
YfM3o3Xezx7TVENXy7Zw+UG2uysV0sPvu75VQf4OZzeJGOI2g4IP7jXrSBxbrevIySpTFyhZ6RYj
YXXssP8uPBpLqbaEEcvX4Gw7OBxWFvaUJQn4Ko31JdDmWgkJnYEQuQCv+GDWnc8jC3g1MbPXgrV/
7zZj0PF1I8sJ6OGtB020lo/HLJ7f0onDEqNQDxnxlJ2llofOhRM7SERnGUgeggYYukT/kMk1iHWM
1QXpbPc+NOZ+2Vk0QcZhQaBWqP0Kp9C1IBwD6osVdAH1IqnfScDlqWOwEw7jRUthjSpzCB8tPDZX
myA+CZBtwlrWlOZunPcTq3d5MEwYTmPF1SahiL5GuebuPX1wwQp49npBytcKjnvvHsjbMbbRKtjd
XCbBCEs8nEmaPHtuR7YUzHuT5T2TCvJVWnbGHPwwBvuCXt47iNo6jFZz5ll5p2rV2e4+VKRuaaQU
IvEoSOXZMTuAipFBw4vXw9vI6zywoLyVX3N/KbtjuC18Jz7O/gvL1vDZKD6ovUu0Qe2LWQpZYI55
mqFAgNIOAvFMmnQwBMlni+ky4vBPsRoUPoPQiOnPN2CACHgVfVJETXq1dSl+ipM88ox4tpecEXmr
uwOHVN0M5xODd8eC1gfGSrw7mfqJB1kJyGs/zI+wTU/aqicnnDPwLKwy8PVrsJFaxbyKT5bNDoqE
Uq5MPKJPhJG8zvrzG0NZ2ak8JxnbCdWWyFzNyQk25l/X0uSSuOrXTpYq2MWbXd/2OA7lt77sW0La
0sja4pI8+F5EsEg8zIjy4YgbdzUGpOeSYkxhgNixcMXKJ7VPdiVp44/jagGKiHwOffhRMVqkh/ME
1WcC8Y/kZ9kmeUwZ3bzIZ7oherwybZiTEgxNAnzIBjOmdtDwEdyqePUFcNpMsjTYi79baH7fFPkN
Hs9bAlLmrND7JPP+xQAFEVvtgLX6iRLcZq4hygGiwfEIPxZ/7/04UNLoWmCxIuTSfldvx43m/bvl
wBIcmtgznWm2lzmAI/gKSCo7rYQO/N61Vs0JKzgjhjkiAGVcAYzH/RyJolx75JlkqUH17T6kSOul
pD0u+Dj/mT3u6MmTvdCyI5tgybEsQptlDK4mTJIkhkpljO5PvFonSPhI+MTXpLzFa7sZ4cq+4s7H
Ifp3OCeliXH4qvZeMQJ0neFEsUYlifA2Wd4G1HbFwVC/khKM6oRpClvF/Cvsnbsc5U8mn9Hu6SCu
DKI4FmQgp75d2MPkQZKiix2jT9wI9rBpDDEKQpbsgfSnVUXa7Yae3w76HxbqCThT5k8RitC95LaJ
vMUdPapKVOQ3fL2jBbg7LPmRUE5zvwzt84D6e/7BkeTCwp7G9WerO20sBJ8fOZFmFPdNGAoJaqtv
QskxAwIS7+/8GDBMR87b7gCZosOj0ooTX49qhkEa/b9HtKsQ/Gkri1vEsZPdntLLHhb7fGxhV1/J
84XREYaGMDOjQ8fkf8rRFKIjuBsri+SN8Tr9loZd+kaSGXO7PHbXdKNwPjnI3UNrOIO9GFLFS/AP
2uoY1gWptJku1Fxc7JtNIyMqFeWMqThguq/T7dIywZAp/pa9/pkl+pZbZthvyrk1bLkvVkTRVnJE
ISCmbSVVRZQaJ/zxhOe9Jn/qszQGkgDj4V3wrSITQXQPhkQ7PeBUijtC8jQxLpFwSHg+ttqdrAdc
hQSsnQSj5rGJXVdU+YNtHJYmIUON2NBlkv+RggnGArVqKXBvAeGYt/dYo83DDH2clhk+Gy2Qhm3i
rLBb8RPIK/WalVV7H0fncaIpEX0rSjJIXsatkMlFKfhGWnd88AtdoYxcRH2CoQgSn3CAoe+05lg7
Re0fSHM4T2UUxZXttNDzFqCcBAc+9XhPQ0SyLTrJwWZ+AFuffQg8SlzOBAikC4WfmIWmgW6sugGP
dybKdPeDPtV7etf2mxg6nNTCzRMwaGHn1t3naPt/47ecLzslRgZqQPqUVnwsCkDy/rnPdnLAhpR6
Bnq+Ft4XlhyX9v62ODff1jF8C6MxJ9QX+rb0h/gydqPKjkizoIgulgT0M9pSRJAp9AwJf/uA2WRi
u5Tmjg29T0mSLZtXVlLjX8t3qsnPufgL56H5DrphnjExL5YnMM6qZSSJxxCEizkASlLFJEJrkmmo
8BNWoZghhYRIRD7PdZ6F8VRp375lnhsbVp5cEV5hgu6DSD7J6J7b5vkMxffdY1vttcbEiRB57Q7A
mwQH/zNbPjOD/SMu1W9Fk0X2HxCgbA0EeKUbYwI3SOOmDZRr8QO1KJTHSY3DMXbW1YHKLxwDb+fv
pO+zfRL3ipBJS15gl93q9qjPqwerl4Y9H/0pzGmPt3SL+fgrSzVmNQtNyNYqm+h/OmxUkplOwzbQ
f6WoGYwMErDJuEYYcIhbNeXcqcjWSL9QT7PEXl/tg2AsFzGl3kyRxhAAFODZMiqaxzTOOklhvw4C
4IohWs1VX0QrP4TXoe7KqGL/2ZnfyF5qTocTaYqmEHs7Ap22DbqehKG3wels6G4iYkVIa2Tny5K8
dv4u7P/pyqKNvnrL7cYuQXSqWg05aqn8qy9UVPzgijCeY5sk87lqhlw5/fB++87M+5J5ggtMY1VI
wqzQcxE3Dck7JET30TIOBAyu7rWq5QqQrs8P67p/hMrisYqfubYdzVGX5UOQjj2z5uaVcSdZ8N4P
LDG5oTMZrE3RpWdL2yYWAzDgNMPEZR8u6WgQmc+fxmpcKAR+r/6cJ3XsCJ9EmyGpa+rIInNBx8Ez
nZEM1OosmP5IkvaDzCY1EaPXBmTTTKMYZBBK4fWs+rPt3Ud8bWYIPslMpM2VPcuaP3ComVoF41n1
O2PmWQXOVOtDW3DWfCz86+B9STHT1LO3CTPPveqEsc+Vpl+rnK6Rtho5pgH88VQgjn4bmfYOvdpK
jKIrr62UlMPAXzGoQ/BRt/FuH4M6XgoqRwE04ylw0VwvKt5KMuC0P0RnWAmZIgC7wRLO26l4oNvu
k2GroU7tL/LKBNISSXIAbO7MFr0v5MS9hylcYzVzox39LF79NEJ8fOsL+j4RBZLdEa/jQY+ETjA6
3cFFhE3USvbym9SFFNbQik0rA6zp7SrAuhpzdiK2OPzkKiBVzgLEMMMZNvUK+WO9SOGNmd9DwygD
xQzXeUSoX2OsS5eVD6t+2cCyadOqqIUFPuGLsC/xRrtaAoG5sig/e/6muJ2nZsYwk0cTyphLcJB1
OFXE6rU0vgMISi+XJHgRAkK3Pmvh80T0wNDf8hECX4vbNVwTPMmXQLyp8zyGUmtu3F/zrBr3R5x1
xlh3xbsEpmdx9C9gfzKuMdXy492Kxk4xTt9FVBcZqMt7GB+zjxEV304UX0i1iTCH883lXop7G0gS
zOocM5lN8nXGOjdU5+U0fEixdqYVZxOpaBAnpPf4d2InCXqeoH7H1l8inLyLrjy6xrHA6ELRvHbh
BIBLyIXRHT0oj6GRzGZBq2LmfWXGZ47UA4omJjuSNW7jC44ErfjalaK4sakwnzHFsZDxex3lqipU
TH/kYmz9biOoTPFlhl5648cfyIhyTz7noolQQfVr3gOiL5zBC8hDZeu5GNd9XBDHFwL6MFlZaTpT
8QWET1nr92wXHD2guLSHlLQNW37duMMx+q86bOwEvxc4DvXln3wP5uyoymucSyfWzch9dnbswPYP
ZRHugSBaBxdBRmJTF9caTRyz8mZsoggjks8mCBhrmGNeqb/bZkC7RyCsSCnQYZ9yv4bz0/jxOUx9
4HhXsYMa8NpZEQkSPk58bVv5/ZvrmNBNerzTvGtaH6pCbjiG52yJmcJVQRp5ehue02jbhLyYFG5+
BBTqwnXO6LWLSS/jN0yNVoOuL7QdWKNHrSMdj6sJEVTU+UTnfGZHYNjtaPJWqcoSWW8FV2OTjoWn
5B7ni+gDtpd3Mlkl0EAzk1rAM1Kq9iQxFJoLUE4Ix4t8kcShWTtU5wQ4HA328aPU5VuOJItfr90s
gUnHyJmyYsUcJawbOMjAXsigRbg91omzvEHP+GHFunpGSETrJiAHv5UxWoEuSJ2mf/8Coka5e/WI
bGKQMs8axA6uy/0vYiLdHFnMDlc5X7LWsRcLAEkuGLQBUq97f8wxXkmKM4gr8QiJuSx5yd+ZVEax
zCrUFe0NKTF3LeGxaScRb0IbrkBqupbRNqS9stxCLNsqoy27MU6hf9VecnJfvKtOneXJk4TKbAZF
9FcyWTy3MDa5yWh3uIWCT/cRXftfJG757JHSiVtQ2kWb//lTxpT/1vehqHrvIP3JxfSGkYeFmlci
2szm4DljlaquBsxR884g2Xf2gNPyA9QAxr2+yxfWgAFul0j/tYSnsqH5JLg3Kh5+WCQ3q9eMOmEq
dApIsKqz2+hLY+XjNJ87/b4T+nmNrdNdTY/Djvui5R9EcDPX83EHlk78YdkECg60q+jBGFPdRqnE
jZgHV/5paH2FFR0sBzRAxLOTSVF1eHLWxj1ukvQr25ODcOxt4zbv9eP0P0TcbO4IjI08Zk7ggdH+
zGyET8bHQoS/gX7GWbm9M1BIAM5Kuyvq4KHZX/j/j0eUmrL5lU0WP+p2b/cif476F2OWrFkjFrwy
FqlTnxDtNdXPUOsJSxO7mmT3qoFmRGy7TdVobZqAcbx/oEs6/bJDZvTU5uG6bJKOfmHxnUPxs0oi
Vm1hyW5c5GsVS2dNZiHiaxhIQYHtOrgloNhUSIr7nAiWuP2XzjtKZw2wVtegWXT7ySk5IV/Piftn
aX0b2bW+crDRYmJiBYCaW3zal8me2IxxfxL0Pr0gyBkElNqsVqJ6oVdP+GRKZn1fvApE/08sg3dB
skF0YqM7RhaUK10vb/gnJwERgHov7EBRKOseSuWOPGQEB6SEEgg1VKZrX37hTBreaGqA//k8E102
2wEDXhYtTSxbYxRkami/H44rWRe1EQ61LJ0vH6JIu3cpecFMLooGAZfWXPDIhVwYUxSwlHQAf8iR
bzjAGIOepjcouigOBPbqNOc5ZuEA8JHPR77LejyX7aWgpXptkN3xKJyNOVtj8HtBQuazN9BnubFX
mjZqcZqYUlx4FIe1w/UFUKvSVAZzSdOgo8CwFcHoT36bt9B/9XFhEdsARxG5pDSnQeMUY5J2exEL
bMWCjamsIeveBzQ8I81S1HgCGMLGOKS5WQ+QVM7Dhzxv8f/paW8tABI56IsjOBmGKHQEwHiGZ3dy
eY4OvexAnhCD03MABgrEqE2DFdzow3A8O71zm1l91Evi/XIpvIAJy4zU8t4h4qQBw7v5bTBSMX4J
nVCoVdfNHsQRWH075K8Lv0IbCPyX8NIashzTpm8FhBKJ0m2OeV0GkGIJuP6OZA8pm93wnVmK4UA2
g2Ory7axFpor55SdS9epFwd+RELYO+zyqHqOPRP9nxvgIGMgap4PIPlFXVdpoaAs6C3e+8AxVYoR
pAIisbDy6TKNNGe761e1J9QDmm4ZRAKk3cs2XNNtpcetEuXZ00IuFNQZqJDVaULpxZSphXwxsUS4
Xk/8fU4vuL2XWae7w9R2ppGlRDMxSkTFL1ssJCLv3J+ozcvVr5dPq990s/KsM0jE83Ljp1goWz2i
UYs6FE9xcuRYimJEBpW3tgqJVsF1M0b++ZteoFjeLcYGZGEjYSlWn+0fm7wama6tSIsykMwUO3sv
4jBNYhIvCH1Iw6bMUXM8oFny75+Wbw/DgWRZ0G37laUOQ9qm9l/OBd81i8mFp4HO8ec/+glw+xX7
O8fEn5AND2usjwLAYFhkC6buDNXZ/apSD33dbKMnBxewiHLEKMM5ppNZ/2BPO3J7qcf4crqcwPgD
rLbGfHIDmQh0VFv0RKPTg+6SEJR2IAz+vZd7cMDifReF54L04CgEISOLa1zbpRo4EHK6o55gjUET
VOr3rbK85f+krVMFNRpXtY37ZC2MYx+OBc+rT5VGB2EUo+aAFanKsllqbraV7OMIZpzmG8uNSgCE
Sz1JDPzfXHwBcA4wMu+bCD872wkTnZjcZnKceCmniLW755XdSBCjWCQzxCTyQWRPnqZhUdJQdlag
ehOfE5tisHUZwzJSWWvK8Lqv9S9jF1NtmTAHaraQNDwTa12vANfOBC/RN1ElIEjE1Upqi9TuszoE
g4QbdM1GKLddJPkH3LEAAuMvra+jtCWQ71s2JfR9TElBUddmt9wFSkEyhhfEBCygjfIFLPF1yL+8
5myIRpLa+V0eNa9XgNcVOyosulCR1FzJobfL0dasSSZwLiVakWwZEPdtDm5pX7Y30o1PErvOk9Am
BBXhN9LGJBLz+x8NNyiQ/543vK1vsbd+Ln+ijq4GVG8LKH5C/g+hqAwtOrUkVQATxH9IsDM3qy/3
BToLyJZojkrUDuBZRiB3lSAlE3zl/xy3JvN7Lapc0nWL/JfS/nf5C4UT8kJNoMQy2L518+VJYHWs
FhmVEyXGaxR7OtKHb2QlfgBA575K+56vW0HKcjGFAHqHBdRusmXyo6yvHdNFgzzirrjsUE8g/2+o
HwPu/YFBes+uxSNOZ8SQ9H3P7NmZ10ATfoNkBYPfZe+VRiWFx7sn0d7x2QETHyq+peB5tKlvCCKv
XOTZJZ78+SFJulGTQ1Rrz2mClmUy5/wW69dzlGZ5sx/wjsILI+2KuNRdapLFTpGy9Hhp5wq00G1g
ekaofg4nIWBpv1pYziKPJWFv6121wbtvrNovuzle51bjEn39wd1VOCuSHwJKsl+pZFtQokeInoWK
IuHaGiNA7fGOj5I1qErtain/o/taXz+rl43YtwxBCIt7/BjvIu6h4d5I42dcNtnBcfQfiCaelalE
/fcb/q6wbihDEIv0en98HHuzGdjD+Ac1bDbbYGk47Oh01b6B6GW4ri9cr8u/wU7ZVQ4UNdNw5qMP
OtnYm062KZyo/SXLw2IoZp2odcyDzM68BFcPFbILwgCMMSnmlEKz/puzMuMHd+nStAlgCo3ntxF1
J9B0BQUIC6KXwNGWV+DBgOHEkNcQwcC/FeLGfHQBZkYh3VjSR3yMvSOFJmJUNTlKYaGsJdN/C6zv
WX2FyE1OMjBPjVOKsTtEx3UkVgMMLanJVA+CBA+ahAx1C1HOi3CZHTiopqtHgAHKy23WYQtt2yQn
CZUShIKewXJkWUFHzVFOeQ3R0bhY77f+AzfLKkgKXZvj+b5JW+Ig/gwTE/CYImrMelSpQ/eVIODf
Vjy8d++Re+vSJXuaccLsiQWrVZ0ogeedv5V/E8cnT7r4Gs05jrt9A7nRPyTX3ou+sqKVwk2RiBbB
CkSO4xqNXSQnGGVItuxTlWqQMP8uZWyxJA+DnReRk4aPNpIiiXxYmgQyBxxosKazxucbD99agHNB
fli97J/UmtpWqiDF9no4Mx/xhKVrfmHQX9ERAmdalj39d/TTBfoBc4tfdm5PafWvnFlrMAAYDdxX
Fccz06/aeyrVJcTZEYsb4vyYEus/d4cXGqM9C5pNE/OwyPNrolnyoTtrgtXlxdENh5o7jseY0TPi
DHTcPDxWwMAvGnLORv3GYX6vS+QAvgbbm+FCNvPfRQnw/aoqxd5q/8s2YkTH/ztkKRtO6g79+aaQ
5qxRHjnKO11Ov+/ImBj4CgUhPRo1FsKMbyaaAqw28qNHoF9D+SHknERfLSQ4D1uj8ey09iXq7Ra7
cVZAtA1ko95kqW2/NHq6MoBfKMf26erLgg5A6DWPshmCRYyamRGiYqBzDTgDaf6FvF93+erGqu58
uWetVSK2mmYJ3dQLWBMNUnwI/17KqL0V9Dir1wiaY+PFcLCmMZx6sEZz93aZO+T2hFwg3bQ5Yc2V
h40Qmu++OG3vgJDtOqG3Ob60OlfpGFfvmK16qINZzzlXV5qwtWyVxy+QHUPT9kWxEfzRrJyn/FL1
STN7k/xCRXVBoOO5GywOlYa6xbT+izzhobqtAour6Mfvk6N8Lp9dZCKaE+tPi1g8F1FnTrzxHYPg
7y3vRJTm8j5+/+AhkGR+Qq55UzyRgpo5rKYBGI8J+grVUbD11psIePuEJgW7tk1HbTj+UBpq7+wN
XAsHmxhS62jieTArlsgveUOU68ccKZHiymD20EHeIcGSNY0vSOYHAGWn3IAKVMHKNFFTWav+vmn/
f6DH610d5sm11mSr+k8DyWyDwku4OognWShXS83S6G/k0PSWb63NV4Sr11sLRvTrlDF/fJfLzl8Q
jRQXjhme46CWX3tlV9iBhqUb4goJct29TD+g4yMsKoGHo1ShXzktKqqSGjkr1iILGpt1GKy/oagA
n4NGZwNES6jGNq82T9bRWnXE/a5W4otYnDnakEr69GUsXWcQ125AJWCtpvHwYVVAvKkgHhYX6PMB
yvEhsRC+9rDevwKOvtfwHh283DGGbysJ2PQYm7go6ExPSMS+2R0oDDJ6kEuEPNhJlmsB/YLmNcVf
1H7cJ6Eojibmndv4cBnGCG2nhi7G4S+1uLb3xrZaxVguhaWyN1JGeLJS7u0a33gI47/LRhBh2xem
jIO5p6dI33nDArA9/21YnED45uvq25aRCALZmqvYxOrZHw2QqUETjiqlhYhSs7z9qoncAb6ty506
B2mjq0pYRdR5UzKmGqU2MmRKez7UORafIfc3iqyhsvvQQUHnkIfVSX/fY8BZ4bGxZzNLLLY/sgZ5
JM3aLB2H6Omua8kjZb3buUsLNERrUJFenq+c0uz8sXWKVKZ/6qAr1IGhW8rGbIFb2QJagAdXDGYE
9liqfqxjFJHMv1F27y2egXDW6jAT8f88+sfTV/feU1YGc2f9CjaBVx1MYCfUQetq8ycfUgiQtyLO
z7KOA2ppkPJ1GMWmPis6NcDLHQHa645fG1n/H9Wetzx+Xt3H0HMEoMmXhbm3SXz9vhFLXYzAUgLC
uko1zAcaT3MyQhPGeFslbSnHW7I+l/gZVlxBQjXrRT5lraeQxKkDppO91Cv9etqlOTtuJXxrYc6y
YNyhyEVTijjnjn+yWkeAYgyuGh+gVCSKcxiwZMCtCPlkonvqT9zfuakP6vTW/KHLcTAKXEXmJeum
jE7ehua46/MVtR3EVtlVRs8NZhUWDHueF9ely1nV7PYupUGQXToPZl2ndDV7ZJfel2p6BGZJf1iB
8ndFjyEc8RVLA7aUtptJjP7jHaGdn09EonsC/CE/nt+O9hJy8f9a2+YzBaB0uNvUBBRWn3+IePEM
GUBCoPIYLFSkWeU9yj05kH8D+9z8E0a83pVqDU5YCfFHhW6lb6y4vibkM88Ig+ChwAxGtMGs2Owz
uaoZm7dRWNbebqRJ9aziGqzGwXK/w2jNM4JqFH1DMB7rQM3Zbd8J7guMNO39BR6VhvNLArVNMf5u
4/N7XJjVF6g3y+Zmau/ilcXCKo2b2fscouiUKdrgpWANBFWNOYFSfl6YraGlWTAGmCZAOLd00hDV
J/kpW9mNvFpIL0E3mzWpf48T4+XD0hxq7mJPSo2DN0gTwNwFPYtFGkQdwGsG1MXCncBBFpiQ0wVt
d08WIhdZKaIc+ehsYwFdIzEBz4morLEuLHdFJOBckzVr8SkTuDAIlhLWBvpJHyQY1ajug+LJGMIO
NKxSqtmsgj1Shj8GdNQ0iaGHZaZbdqGcowxEpUAScvDgblTs1H5V2A2jEjf/SM9skrKWU8oHvU+J
aI6TWmZORy9862WvKUDgiyMqco4aKGaMAr/OsQSLrmLkq6MgTJPdYpdkLswLdFP1JKBIdU7WJu3q
TJjbrFmwNfmyrbwGRp3YAoF2/VjR/MPtwl+s3ZRbUo2W/XyqNOKzM6oJKQrQSz45E1zXfNFxHSBO
EVH+a8ItD9AntK6BIJiex5Jb0L8vFmzE4LKYdkq9YEjfpNbXZ3K2KyZWNaYSxY+HpN28m+Z2T19N
ik/7HD435XKLqVtpOQIkPlzAgP41JzO5NQj+76/NyStC3w8Yboa7c5q6JwunDr2l8tjI9VLap+yq
K+s4+kyKkdZ+2B8i14fViQMh0gU4S2mcsjlcuS08JJHMI2pVrkdVzJx4jcG1QEms9Nvicn8NIfsj
ULxfIaELvHpGA+qfTPCM/hC9sMPJ1fVb1xi6Onwj7mH6YhJbSiR1I0DbLqEtDf0QAGAzpmKScwTD
oUD3Od9M6aPi5BV6JFBICQbRhJbqQdwUc7oFzdJJTJRGb4gxKI7CfPu+wM4BJ3TBWDoB5SR3HVle
9XFE3NreVGPGI+NKJ5NwtBtJl+LL81x7qO0kWwsDlyl6FNM8ednORDyti0q89nODfNB/Eap4CUHC
inuzQu+Sehwvc+Ngv/rows3+YUYQVYD7HjqW+K++/0QUxE2QTHFEP4tALYGMuCEUXu1Fijmd1J/O
l2WVe2UWGXm2JjQfLaIb+Ph0t8qoiMtzjxpjllhXOCsPs2ACOlu3VAEYFsoPG/TZz24ClrjCqQM1
85S2qbDyOk51mr951szacq7MAR8EmFWfM9dQt8dqcNVCv6B8E9+1ymd66RcizNtmx1fVrANdLsIi
AHtW1RbcK/8hJnKKt1fYFxyhg2ivyNA+gUBtO2xF9xxwi6dhEM5ZtIYQaqWamg0dOxQOWRly0MXo
Cz0MwZ32IlFcSoC8FMz/Z2kIrZmW6PGlrex3v0jC5z/Ucg3N4oV9icoFxaGfWa0waCDcsQjsfjXg
oxFM7ddMfoTz0lY+m2FGylKkebTSMOy9MCxhHmcBtXoUJK65v7qOS6voXSAWMemtSRH6IbgmiNix
QKDgRnFkTYlyfoVAHvHaB8IfZ8KXVcfTd/8boe5+BT8fbAs1fjMm4BYn01vVARiiFLKoygtcxzKh
CD5uQ2CfPrHmwuPgLL1pXhhNmpEfLrYQCb67u3quCNVGUYds5ktNA/3+s8md/oQOy509CJVVjq+y
4C2aMzBBTQzTm2qhWfhcHcWdHkVqRBixCnXKchanI7BiYY3QkHBhW3Cl+386jrfwbHdFkOXkOaDm
o0yggdr2oC/N4pLBugSUKdxTdneCalTER/0NM8KcUtzexIAtNrSRWGjhKTEVZ5qcDDUU9fRJDvBf
SV/Rah57XSfKS50oeO5Lhd1mCtAHB7cwXgQ4v2BOgYpD7Y3oJh0gG7Fr23gB/rTTzhgqYYbKnfeV
2HKOmZWLIJ9p6xzx3vUGxzfpjPeNZMg6vzbOudx/akQGY+T+TbCJbXScAe9Xl5UNowrUD/6Zczhr
yOmjaw8nSLxZGtK1APlsJAOhVq3Vxuf3L5Bmc6tOd7l1ejFMkiTP3UJblkrtiUjQ2rVJyIQtxs8S
/HP/Dz1X5yVgGCSmwDMBBlVyttLoYAqbaFYdKm1vs5pU0BT2yJHQIptVxBM4MqmkgVL73M/Vb3aK
Uju5UdThDElF8AAnxkbInmMYdqwRn2j0N0sjCBSnOdUhNyKn6RaLzoKwZVLO/vtLmlGkO+PNJjc+
CbqoaGEYtQ40lZlQUxtsYuXWVwLktgS22oe1CHgvTBSDFHwxuJ+n0SLXzmDIFFEU4GghZtOAtBH1
O9BO/nUB5IilZihPrKQHri9s2+c2HKMpjvFJLfVDsZvCxSF7RIw51/ui7kMW0q7oWfC9ioayuZhq
wB6NSQ/2EvD2PzEKcIAIMWyXxVp173zoWnQbOGjubJ9YlcrGNdNKJkz3Q06fZ+Nm6DTK0+A0aOcd
ARgKau+BsoNkFGDoKOrBkoS7TKhnLjqhIs1Ezt0miZHedOrcXDoEnl8y+UCUwaqKNFXbuzvhb+Kb
oNtpBzBmcL0He5ANXhHbPq+pI5ljukzbI+AFx3jhXg0jXWvRv6WusJRnJX7fO+Q5A3DnpDh9GpoS
dl9vfYgNW7fgORsiijhp5R3s4VXkhq3U5qRY+QAwKLi56+C1hpEFM94exTBf/enMhq+Vg8b+bHmK
g9sEtHywACve1cOVd5HHd5i6yLXx3u3D5NWYIju7fUZPHJLbIDekQ7uTG4LewvSm0BzJWzPyuE2F
yrkKYw4CqL84gMPUpcM/KoGVpp8Uvgj6ubZKQsinMVh4x37+G1ND2E5h6cpbYHWQSATAsD3bcYJ6
SjrpgDm6biinhIhvjRCYhmDRbyNf61UVMDrfbVOkvpE8KlZYeKXtjdgWm9vh7bcXguP5k6a3+LTu
UENiMrvvDoh1MkX7wnaIDMK3cbWyYNcLCLLlNjVbqaXe/lTtfhlL28U3Jo3+lTp4Lp86aacGo9dq
TftDxPdji7liGTwnkPA0LUSeoLV1UToYB00A8QEm+PDcMyS85Mdf2cBEQv8HlOJ+YWKQKod+2RAe
qbXEIPqZKYY567eq6OpPNIKB+4D8tssSj+aHmm8LB5p0MtIbBwhzdh3IaUzrtY3whJ7hs1uaP/yn
h999ZYcTINJdI9tdw3LOOMu+hFFwfMm+JfvoRzMuY/oInIQZK7HpQH7X5L9qplMHiw9RSZZODRre
cDfsyljQ1eXB28PX3W8T61v+pncpKgcrtpn/ztoo2qf3cyhDQfauaFoU7Cl/qa4k+jZsTcnGMEAt
4Z6nODsvmk735Ehqf6yDoYm9QZWmJUT6SONAK3USA7xEvToQbJdJhnk7j1FxLUtq9oqaRAN+KSph
ezSesiXFLFl5QuUKN+56jWYJ9n1FG7JjEalU2RJmPDHsrFPWBeueSmXcTnM4z3oF2fic2BmE0bNa
Lp176C4Y2eePmLmFxebfWNKEq/Dta56ZZtUaZ/E2bndzBHbRa9ALYv/O0vwdtNU5TJSodYRLh5fy
q2wuyssY1179l8iAL6iUmOg8gVyqvXEXaab1HwzRvCeNJFxGENKfx/zrJ2q60Yu67X6QRv+3xIUy
8ywYiwBiSgKdEQBphyDw8bAupiTh2/5k+VEYs7DMFSrCW3nTwrbAbERu7YHI2kAi8a79ZfPW/bpi
xZE2yjzlhTI8g3nv+TZS/6pqDVIeeO3Flw4d+E2NYQUE5u855FtxoDTUXZd8ykG69EQQ7kvP7Gbf
B9zo8cYPSC32Wwwgf4ZJ3zzq04y4238mnd4CZVMrLINajupGIyZv/D+ZaBz6InqBpc/VXCzlpHb/
twN1ywqtJNYD0M4nwOIauKjinNfUnId4Al6oyVcVWLOXi9J9aQkPqtzub92AeRJReinwEn0utgD5
/V49CSBRVNhvTeaQciGB2W0rJu5RwCoKam/kTvIUFTJ+Ytw9SomRpdrJEB45S+BUaH88cSfZZXqc
K17aCpdNIJ/OlXvUQd9vnECBNBQbD00vlyn93bUwvs0VbtW+UxIAWUSJthMB6SjyrL79R8aSPeGO
WNjo+llXSajoMV3r3Su18O4XDBp0KDCHr9k5jBm6DDkkmjyJtU7pZoNjs14QaijCrUBDVdVOEnZu
azayJAPa12w1uhLlqbHqrda6l35ro6whi5TLcFiGkZW17iJnM07rKqaxSTQM+PPgE9tGXUKJqqHu
K9kYCy8GXX1Xx+bhzyp2BHT2xZHS1irUGH3v1c6YWxt3BQRE7uIvH4vgFdOjUltBz2v3xJoE577X
T0BRMlFQ9aa/IQ+RRDBW6fpcaPxsZZGiPU6yl8b/Sj/UVPo4jW6rJ3ZjlG6xrap3vfyZuaEpIb5N
pH9jenmu7c4PNzypZhUQ1ZW5Za3koEmu8QE0Z7sc/wwN+cJJlBXi2GfJGoxR6Hf6/A/WH1msFb89
YtAU3m9nyvEkq6qpeglCpGldmVpo0nFbDeRhkVVJWuRqVfJIrzDIeUTDuuoOrSTk1Y62SjJtoqY5
b9No8ELNd9T+ys82/5EWTSD3gJeCIZx0WR4gUkuf9Rjc3UoyzSFkFuF9zZGu1TxsTkXRT2eOXADD
33AXJuGruvautoGbm/cUis4SdBDqh7vmyP79NpHP+FLm3geuUFrA/igfhcJySZg3ysVaYiOk8XKr
4yr7pEaoX50eKZ98H1BJSRgKoLae61QHwxEb8sLn48WYgkVtPgxsl4b+QiblpK4GHNLqsgwPxN+E
TvRGiA4k2ubke6UXr2QYaMTgRARo5cguCHgKakxnCLl+KB3eSKrJObkn/kZKxWXmnpb8UPc5J9qi
yeG4gdlXiCo0uws9l3NlfAE9IheQ7VdjsWoyOeMuLs2JmeFASczmG+Tj5Hww4wEDChaxLPZ4BHTg
rvC80axurcZxGKyY7KdSXpcFENQnKj53TlV38njV/0h9oO3J4ymLFosqBTSS8MdRKvzEi26Oj/o9
6IFY4f/k33NOTM/gIZU/qcfmPMG4H45oSr/IcKuSNliglTQoblw++zVmx0LHEJFvaProL4+9WQ2X
DrTe7qIKgUQIitpL6CDTLieePOrlLsRT04AKIhg6sQ4S78gFnRHSEsv9xytD7JZ/rxwUdN2mw2xJ
0NIsq7C/C0mT/BclXaO7SeRlUEVaYm4L5ez5FtR4H2hmdk1Q2Ag82fsEqS8LzAOFwYXyeMFIi3Qq
Woror2Bjs6wLdMzDtn0S/sA0AoW1yJZ24VnqP6u8O2t9ebO6ZXMWrWWTabXkR0KKcNnvPKiqsVub
H6om3p7vFhyf/eQlr4ThrkQyWECLvuHQeRoUF0JOGtx8m6Dvk97UxO9cPUAra7Xe9I9rQSF1tLNq
wzKG6S8//yz4Fm9OJv3m9HzIPkUyAtoZ4OVjEBpGRJShcEasSpfbkhzGJaabwHILRqWnVrqjaLwG
2wXKAuR60gje1ENqt1/dMt4JBH2JuquqG1IrVjbPAghlmqzXYoVTZqI9HRn2CZAh4XTX5fn1Pdm6
Wf/HvUVEWNXvaXMKCLsfh75XdkPq+5ZDw9NauXWUzJISaC2FaSH+OAEXNql5OH7TyWMXR3FRvHrU
WdjNhjd2S2a2G9TZdT/43WNz90gXC3iRI8ua71TrLqW3UaDmWWwGxUQVbYWT3P7nvzhQnGJ9BxPV
u2/OWR3ug7RZ0IxKU+RioLHLYBZeg8m097H/YNVqU+nvXHxx+8cuc88cmly/G7FtPe7Fx8NGxzqo
82pNeEA02lD3hEX2W/kAriX2TxlidLL4uFbZC9Jb9DTpD0yYI4eznEdLhqNqC7P9GddTfocxSAXc
zrPRAbym/IlVEiLe67ItqZf3t4QydSbvjRMd5xaNiUwowMKDnxiJOhB1FDwNMPCRtHB5vhZ9Lnzh
1lniGDL+zX+yZ5LdIt0137XwgXksapPq8JXnk0zggt6IJlxq1TzHyu9CR8sjcgYlJqArehgIypES
YvahCmUd2LoHqtoqT7fyJRHGNtnsYFk3hiJTwLNTKuSyo9HpMQBeQZq+Dx5vc/dHRG2R1G9Xaahf
l5kK1olnbHniHxIMK5X0upyiw8FtpbaEweitpCxPirJQOLeQuPp3ABo43XWcXsIKoVf137LweGhc
1RVrXatZJylSyygmXDvDQiNvdiiyoqfY9HfhT6M/2WxSG289GDDbmlNLaP2rd2Tcul4Esa8/yGL1
bSqZ5XJXy7vi5ue4oJZoPID0Faea9KRU5tfVquE4wzGsbEUG+vltPj2/KQEf+MQlTLsYx9KHNJIE
bEXhi993gttpwRWvAcsYMY8FCF7YRlCLR+oTsmxRSqW3ic2xRzRH9h981iVo6x1RgFC/r5UZ/oP1
zDFNYJmnen02kDZWWmCh8IsFk4IGNodvHaUR4mTRY3h3DT6/YIVsqdT6oU4vOqpGPodbafwU9nNC
LHjGS708i3IvR6VUEeryrf+1n55AoCisCHM65eqf1e11+2o/Gq2/lzTtvglUwj2sXuwfpuwT/CgF
c/rdzYOr7ERlZZQQ7S2/0lh4WX6CHExZ3ZZYYKO6bJOW+L12cPto4fI66kjKm6V1cL0GqLFO1oFZ
UanhgUdQBFNnM3QxsetTgq2cuwU0IeFEmDz3LutYlFpw4jeXhst484ROEUDSo1jOqA+LWgnCTwYS
XD+n6qmE77+wpdjIVBM3yUHUSTDybYxmWVBHv8XmXljtD8TktWH9aZECiuc3eATP+bx21Fjg3hgH
3l1/bdyqnV5BgIDcavZ1ZTHkFOlV/esCMUhogEnbDK2d/rnXFei5/DQo1fLt5adcXw25ujU96cM4
LTqGlbrpJ6/f+UIzgOdhlu9bqBv7vDvrzn2T/G+9UrmUqlZ3yDZIOCtc/KMSaaLkCBtdC4Qkdboq
u8FAzgwjjs51jhCs9tYrFA2dhKZbEzTOOsvqfpqp/iPdnB8/i/dyNwa5DEm6Y/mOF6EXrztzW5b/
MvxYWmMyfX4QmUM0NZAn5GatZl7rV8O3bmPWDjm0NUmw4xaWDPHYwPWT+GpW3l7HN2E5zZZf/1XU
MNdIKbe59CA7zirSWKnPTn7s+KKdJ9XghQvajfWWCas45WmVhLBmkKzLrNVQLYw19D3AyZCh28hG
1nI3/7ldQeJXvABCuhdO7YaWAkEfzPXXYgkLdSNPCDc9igawoHYGJsAH0lq2U6zLHo3G/t30rhmE
MKPAfoecDAvCai0c65HZ8KLVj846aZ0dz7hAhvjpbKcr7A4EzF3TYQFrthEqavZEniJOcojP538R
S4ugLcmk36E/mINvCwIHd2E9M51isaqKezTVu7RfCBwXHEd/OTFG4hTD1nImrkzSMDXRC4vgWokH
J4lWy/YsFivuv/Dg24r/roiGBYOC4cYV+N/UvvAsIk0DQD3sK7ZCurB4RsbC2ZjVtZWXRitP2Dds
DRcCLdvcdYwxziZYxfyhNJQ6LsvM8nTgdNlG0gWoaM/jc/2IMIcT+ymhsXgPCURMaTckgXWgb7sU
i8zu3MbbUVUgOU4Ih5M1FuZKtvoOoSu+7eV9fh6yYr6ZcLW88eJlubTbfWF6N8pGitdudHDYME0H
46HsKYnkF3Vy9A4qFZ/r3kvh3UBFVyosEn9BniVcmd7QR7UuiFQ8/qocWFUX6GJDFZfnA1rWagcQ
MVfX+YYYYf6BMHjrx+xIL3dzeVS1mnNof+1KbapzxQhIkcos2YryS0xOBUZ1tRCQdtZWVpYg74go
Wpp8X/0va1iA+muSsaH1vGQ6kEfLmR/UL0E43ofFvseqe9DsDkwXp+2QLP8ciQXyfbL8nDYUJS+B
NcSs3oUtLeNM9aunYfCh187DxxaoQFU6l5hL2iHltJAoSZaye4ooL1pzu7b89Faipbaa9J+hCtdh
UrL/S4TUtaI4q5bx+fz3MaAtslkbAdJoi6rFY9dp1UTFAYngsZuFwvBK5ZxOcRQogkF41O9abq3M
IXyMCqZb132IcZFQtbRHm+PlsXePrCINhUWWOzfFBTDMpyc+gN3WU3c+s46OOUKmNhUo5KMq/fQK
iGw1Efq7Vgncy6fWN/qGOdRVdUfZnZ9F9CXtmNyrpc2xFX4+eJY6fJJAkWLYbiFhJzZiwVEPSke7
JVavVoger1jhfZDpAbzaL8oOgI8zwt4cctE5f9WceRI2/VbJvpzdSk+za4GcfXtDAiIYxbCaQ/Oc
EVnRZH4EsA6p22aAM0QsYcHcjR4RUKJPE4mbkbJlfca27/O/a8iYF3h/wg5LAr8hj+JnzKVSFWCd
tQDqfFC8Qqros3wvBGMabRTe1jsSaIfOqmtmrY8CksiqCcVDHmee9I5h7FADjhTDM55qgELyi+Il
bZ1a9VTZ4UV1fVrYBSw/t9tqoloHmXt9+Zz7cDumqFQeU5ysyWq/8x+kXjJ74yOg60ZELz0Xoj0N
2xIRn89z2DW8vF5gi2sKQdDXkSNUVy+AVJAw6FgFVePoa0DzXd0+79MgAkgA/7CI9S8vfss9VN88
NBYC3ugVnZE1xT8KZB0j+V+BFCKhYa4/jeePybieqyYJI/xioDkmk+PcXv2XDVGFssypou8fTTgY
8UZTYS22ZbZP8koObJD26hyr0uGxCssLhaJLDId+Sg67zo/PZD3MPQBF82KY7lea39bx1/+qAOPy
cpXUKHU8VrCFKMzeXk6BCj6lOSLDCU0asB4xMg7SYb1MxZqCV7n7RK+yRpfnDuzzA46+Gu1HrL+/
gFQPfMn+pO/qeu+qlJmTlg6js/BgNg9dclnmXNi82hSZcKg4YR2jlPCs8d7oJWHDJ7r2x0HemwMx
E/O0H5u2yFsdfb00q+lknuc0Gr1KP1dnmpGtOXwZ7psLN8oBzUpvXEA1nU+lTQUH2Dckx2Ct8te7
gDryJcH4bBBa6Ke3VpDK4kGbnohuEA7keQjp71GADRalSVX/C4Z/LzzwX2ZZx7RM3xsQqsH/82ZR
UQ8SbKfrReQ8WzaPD4RTwcIybCH7dlrvBosLtmZlVtWatQKTu1ImuSzCNImvQWM+GyjNxf93DjPa
EjF4+dbl0hoaoAgnMFeAwQ4sUxMadAGS19gmlBl65kPfRKwI/+KiIPgGz9L+YMbDKjT+z7+0azsV
VfQd0nAs8EHt5wdGW193bVfmyXzYmb1oaY1QbC6WaB0QclXjtzUv6wqkVrzfFzYSSbkfyT1EU5es
AYiaeCQS5IvbK/eIZ6v5K5GU6s4uH3kV9PYcJ6BCLmXck5OhRVj1uavG2Xeh1P+YE2Cs0O6Rb9Fc
s4qQkIsauvQRsukBq96r2CUjgqqg985Zt4tq+YEk1wRTYqm2+sztIirgumeC5MZH7Lmzjf911gFO
orwqlshDSK4x4fwq+fHvMKcEBLgI+lUSg4czZudWAZn4oitMp0nyic9qU9m0votW6dLAOwdCzxoC
gBUuxmbncYsz9ENK48Ph9DJUJyeqvsXdwuVE15PjNVRRFqz/unBSNl9wMgjS4QN4uNw6HWGQT4IM
imY+ti+1qjS6TQHarTr5pnyTui5+OwOFNsdx3LilKfZbPZdOM5K0eBimeMjHSWxo9WsygwXmXzIb
bp+LIPJlEiIzJ3lAPG++LC/Joh1FzclFJhi/tvcqGNO+RANGEwQxKZreh5DVwcYBAM80T1PTmfTp
p8cQanQVddR1qg+PzdSuWM4bWUouA4W7V14C5Ob/QmfhmnjlAPimEJ1NRLhqTMAmNBeYby1zQuAZ
2V6H/t8t5biaVcnHLCAdyVS0sImcfXFwBXCnSMszvLTrSSTWuCgdw+HSQ/6EOlcA4tdSCDExIcDX
HlvQmeTj+vMW+VH/+YuRKWOem8uAQ03bQhp3DhRmyGEbMrSEn2j+KXQRf+KTQnS/8nlGwFL2r5H7
li0BGFnLbCXrbNVEf2DaZMYkQVyaLDtfl88EJcpYJBAgvYAGqDQ4Gz1np0JbQmqSfqG+CnvrpfR4
sIhf4AgjV9AHasrIVjQybkdfkYt06YS0ptg4up61ogwvZ4Q8DuToSHGosumS6qPorbdfWf1nR9AM
jYVRPo5EBnygB1qBGHbcnukOnwtOcSSE4Ea8CsilCRGWRIYG5pVBpjOytvo4guZQg7/O/rP+tX4n
r/byXjni7XrQPXbYqlKZXkAQo4yiIfsXuMcFGDhwE58SXM2MxEQwE+KUT93J5566QYfF0K4Xizqm
tguUqEnqiHc0NctwBgk2fhmnbdXOG6LtY0OJfWGAuZqkXnWUo3mLEf1WOVLL0LjG2kQPqMXYQiR6
Q7t+zusxqJU5ULmt/XyiNhzNBYyCIqKkM61Ru9zO12Hx0SiwY71zZ0Yp/kDboPvSgTMX+p2NDzZQ
RyGrkEcAkK5SAYKtxaiiw4s5CNPwyOoQaDDu3K4EdMHL7jsjviqttlqlUdtbM7CFEPKg53C2cH1B
QtExRkk1vv/52Uc8ZVD0RYQQVawmqbiKZ3utKRna+SqBYJz6U5UiC6DUFkxb7W4UzaGSiw/ZfK2c
xZLHb8nL8Efhh57tYmrLg8Tzd9WAc0/w9K3fny/0LbtKqddHw0w9YcHos7MuT5GFAQkwiAwbOmFA
Xjkmqp8FiDvm3+kY08K1JKMyMydoyOHVLK4dBauZir/Tx7EPO6Ru3TM/2TpSQWcIQrmw+ApaJx6S
J1ak1nNqBv8TS/ekL6zsXdOW3lmn1QnbQ8ncT/TM7QzAr6lMOUQmyZY5MPeg+Bi6uLnxc/vshaBL
8nN6kNvcrODFJK2miA/GVSfd1PZkWlV1r08tYrEwlKZU2CGeqxLNYiwrJ6J/c6HSQ3jIlWSgaGDq
T4uFXjIzm9nNXa/B1wloCSf2E5v6cT6ptvcGuKvC+IVkgOg8jZHOfQINTulLOkDqtWJeeDhI+EDK
49/ldBVA6v6oEaBwx1K3PRTs4xD9UQ8C6csQkLgzCKcB5zfXkBOB1/RvyA0PZgCFK0Gcg8NWsj+d
X2qxgIjATNvtU653CUuol4KhpR4cmGqlfE9/v8+oIaUh/coI8GBBQzymr1DtCWjkVDE0iKbvus1u
9qIJih/1fPJ5lALbgYEiIFb/pVOW31QxfhrokfD6t5I4BI+Boh5Ra435ym9iqHlZ7o/umQtaA6P2
IFt4d+MAQK2hbOjVn3cDycWYTMdOH52F0mTmF+chB2X/QuP0jTOA1SbhgxWk8zJoIO+TqVddklkA
fBJtgjvj9EFWBBK724X4XLN3CUNheEqiwbtmr7DRfslhMMw8rfBghUKoAlc3UitcVwhoW0bfbHTU
lmcOU0HG4ebtjxNB6KgWjnPEeDi2qo1qbNf/HNO0KJrc+RgF98hrgZPwVJhJjWk/b8k41MoFuea+
YDVKYEdRWnv22SqYI5Jo8Yp0pCdQ8mSQWcsClXB7zJNFrIoYJX8SYJ8pjMBrOa/6R8enWhOETkfW
kfZItLQQu1q4xS9EyO4c473yso8DmTjazJmFqcSGNp87LfhBx1eNX9DM2V1QO7Rp+1iglO/sV2ie
dwggy30oHUUq1KDCNLvdFRhQPuZ6aUk6vuAT0lFIwx43OhTZAOkj8/pk+sw8Cm+zqmqZaaz2fv+v
Ao3UdXjCrpZQoF/ELZU+512n24EkD93/bJ+kvrJgUmKggTzr3cglUwD6jQZ+6ZwsisFLfot9rLHr
hZ7zBXn3wQJlnBA/mnu6BEjkqcXF2Wy11J4oqVRxz4FTwdre3eV7SZiNlYc5yHVQFqEpeKGPlz5p
kU+iEeZ6DD3/An3eGXSgDk+WDm7Q7qko4y9tQ3Ke3ZQGVIwAfyEYkM+5d3QQnJTuDJjLNd3/Kzl1
+oVYyOmtHI1PfIVnwVyT6VoBsILL0Qa2VCD2nuUlcv0o3WkfXIeUnQYUXohSxN/XzCFfYrN2t0r+
WMnLyv6akCouH9n3D5OGU4I8ZYQwaV9RXKWRCqX5ArYh/26ZcMUIjBHXk0ihNiDmw+NSShb2/qds
OGngg4viWHX2FzjdeGXBt1hNEb3flfaj0lKky1IpnG/c5GwZG0IhNw3i4sfi1PcBigVccC20oe4a
MgkUKiAmqLzGX4nZd2DJ0audm4Bu0CSBDchOMuTtVVoXBb9+9/Ql/1vnV3W3kfziURa5Jbd4kQLC
7bdSum9qxCb0d0LMVDmSZx8/yAlbmrQQPt9UasUBAOhn3uGvwpQNTknS6hSSYzM3rac/+ZZiFlx8
lSnnnH+MPInRZ80s3VWhwGSMS5LHYLxnFJYNcbFdz040nEBpsYijpnwyrmxK2yt7B5GVfDisRHSb
aMypwuyoLHxb1mEFSL2donAB3/RQ8UufSy7VkPJlg+/RxrSKmE1q5TTkhWuZ32ZWAtfLrdfc8D34
wikbyZasbYC8c/xkTzWA43Q8PCB+GghKEwL6c6dswBNyOxVoFo5zFyHBw1SpPCmYB8KIi3KcCi6Q
4M8YU3GASXkz/+INk2P9nbZ1VCn+HK/gakZocF77NYtyhIn4+UnYFizmYga1gQvYLMBEggc6qXal
cDGhOASVDS8peE1L/p+hVYjwkV0gW7zaGHqP0GUHc01wC1mZFnaMkQFkNXGOzwT1vsv8i90pM+aL
a+6mmYBkAwILwfgJLXIEfLVqxGJKIrIZXk90JYXV5W2pyLufhSWjudgbomH+qYz1eMC8WVKTDBE9
1ZcTHXkFZqA9drOA60a+CV7KY0PQulZ4wbR6OpuotTZxxbcd7EGsyUDBjNuoa82qAQ28gKdJDTYv
+ooeQE3J4XJfYnzKz8mJjBQNt9UwTzL1x53rNglX15hvrsWnRcmCLCc6EoxFHScaqnfpolSaipUj
3BjtHwkU53/4y1fGIAvhvYxPv/YMHtvFS2VOctob/sNnSpSwZhom6RV9P/tETZW6QYdpi2yItjSk
waGEjdidP3s7NAeSj/IfXxguOYhPIgy6RV/aAm7yVzdnwvnKwbvql5a4i/i+KGMid+zK7dpt3pk6
FXt2mwaeCUK8F7EPNG+/cU888yaWqIjkV9XM5Q7z2gsklPulaN6hUUSIun+jtgy/Fpo8mfNvaAea
hTZIAVdu+E+O1CbZ1TLCtP+Zd2VvYrN3NNMeoS3WmZaJ8xmlWhu9pvfuyJv/GzWiL1Eg5XANufPj
9QQ0owerrzOM9LaNG5Mgc+dhRts4YLnpmiyDlqk4k1YaOd5iPlvm/6UrTtIZL22eBoIE1p2U7LM+
ASNLrXVU0UB9c0LOrF4MnNcycdNGFIlOImi6ZLbEd1KMfrXhOBJYEGAuK/M4ehnVpgHzPj9pNqdi
DNLEV2gy3J8pwwUm6/HwDBZwtjqguCBqP8oZaCa0mn0mN5cvzF54WeTQGyzhkhgfFlq5XflYzPC/
bIvJ0V3KorKjWhjS2LCi+ez3t+kEfIUNRSyS3FCsqfJDM48jdcQmlp1Y9+avONN6x0otu5sfq7QU
fx+2HEVWtnLr8A34aDSUcnO9w/Xu2ZPwOZWaNEFygCrkz737FzNLJOZCon0Re+FxAGLcqLnsQxSa
Nxg3SSD5BA9+DsydA1nu/XcwO5/TgaWnatj11su6CKD4kTvdHXqlVwl3JtXJSANSzRSCZFJXPJ1/
/Q9ENKGpnMpnWJAe6iO0Bm2ePnyabHrIG5pbZKorKTtc3lcnf3xBYFTRm6U6u7AvKkAKCqadgMSw
zm2Rud1iHhdMryuPy5MRXMi+xR4Vf8OGfoDI7EngPtQG9kQczeyqYtwSnuoql8CtXhoruW/BAPYX
1Kieeirtjq2lUH32PNo9XbgXdlrwZHe7py/4490hfn08IrK9CyDQ+3CVV1A+Xr/QrZYL2NcEg/sE
32pH6RXZcOW/1Fx0Ho3d5KJPeVoJACRTEjp8R5sdRARzxF74WKIqUE2KM3hKINkwrqWAsdLc7yUB
zK1VvFseRpimtTtCYCNry78xqYWAWBDM5or32ozpriIzwbxvacQwtL9qhDtFuHpxKdLbIkVcVNjB
SC/bsyT5riFrVixesjLNP7kkNivi1eW8NXe9euiy9hExj4pXHui1h5cKhCFVUoNye9qhjGB8Rfdt
Tob8lwQ1bjsD0Ftdzq44mwzmIRsBkUjT7jRtMbKEAWuQCf/UkWSSn8Jq3dOGG5S3xYROQVsty/pP
Hzj+9wylFDmZtRaQAj7DmZItVw3l2EBnChzZXKTMEahSj6culCGZHnJysJNtPDwn4RZUwNSgSwN+
Ko9de/rUJplwDrqhmY+sWL6RkjhXTR9u8e7GBhD1DvuIr/HI0qg20NUmt2Cks5+MitmmKgZUA2cC
uitqAWAMYPwNaFy1dZ7wGidC9Z/6xSaRQ4Lg7WDE71M6DgNYUZqQf4X6LkPWtJ/XYTzjEdWMOirR
W+F1sAbcz8c9pqDDVs3kV7HPliwujdd6reskNLHHi1UzzRLfrp/7W22rVk7WWkjCMN8ZjnIT/iWF
OY4KH/BWk6hJVoDt75UOIeKH/zwTS74Ex5Rv7oZOOHqJIZ9dJdIATuPtnDZuozdhpAfM3DtVHebx
RObG+xVtjGhui5flKtEfF1AIQrWZhxDaDftxS9OK4lCrpXW8QzbfIDCuFufVf5vy4ELPfdj+d+kr
zxcUX/47enJ46kHkgJhr3LwxWhu0U2ok5kiHUt3w+7KQLzM9kpn560YhrGGrIZR7/n41lB7RqKZQ
PobgP2oVwEWUboSLgNt1qoxyzI9RPyRuS9yUB4cs4GIOPerxsUYbRzIZ5dmaBRHnBTlyDFkrTVVg
yxgWKbx0V29K/6twNKVx9k0EdL0pdOrNFTx4Ql632acJrFjkKwXaFyrZOwjjtF51DKB00IEJxFg5
AdTeYt8IF4Jz3XsC5ImL0mTawOQsubl2FaSN3UA4BIRknCj9XkzOzAE9QHAaNcFDUJuc5m0u+FED
APpgfO1hDtWubvUGUyOAZv7ybzJhNCVkY0z36BPhSqI8/ZR2awJuZfCYyAxetMOnzymtAAa/4fLI
Ev+1YjL917kM+QBP3mRm7+OsixjtViaE9Jazk59aaeemiCByyT53J5m73Q9zHPzzr6c2BEZDGL1/
RbBdpzderFnYFtvK0jmnreMODuqqiVVSOJZKAf42ATzC3QfTBu3pbEws7zXFSPhow6VzMqgLC5qP
AkUvzTNB6ieJQ+wMxr7PL2Lj6xLp4sJY4af4VMSVxjmVaJlO7OIM8J/sDPETgzOUfqCHMt8aRL/2
uYcI4QWqV0kXrYWkrUg9bllZerS9zRcHzHtuPek8F0SSRl774/p3X+DtvEwNq/Fx2OkXUn/pJhwF
D+2gn9Soo/zUp+BkfCAVFyB2I7X44XjtiGrWUolekfVJtgjmgJBiltuTkcG1G7PBRHJNHbVWlMUi
nTChoMVTwuT9qv5omq9PqojvBwWsMg+wmbQthMLNUUOPZ8ayhoNc2M1Mw3DWerznysnzKoCp+R++
/zt3xYrfwefpgdRgxSnyx0RryWI6/Ndkx0JhGCrUaLC2TVClp9nQa4kiCYpQPD2jhP3e3w/MEhqD
lIEUzSwk21wWdGrg0yO98fOrX/YSgFS5PFd4lx1yX6JCLyYO046RtMHzQPiDgfmh3OJLH5cscKks
FEUAZyzr/hPuzGTbAjqmT4goChMguy5/TjI0q+UztH5eVxCJydw1PFeCRCUuBWmjkYrwmg1/1wm8
xFrdoA86skKoRZb+WEDUm8OUxlHLHrPq/SQfHTpsRM2X6lnrt0QCFCyq6BQ9KWJQRg6kvdWxI9c+
sXfNOWUQVrt3iYwXfT/Uj91CplaOgMUmayDod8Fh98mIAGBGXMVhpwbnrgIur8jffnSVKgk9YdyR
YW5WJv7p8AjO5NoxKGwXYdznkr8JMlj87KToPG5ahdryrPQvi8gIqBnAR/lt7Z4uXSP3tL7IwmW+
XXrusofACOKXn3R5l4CRbJy3QFOIXkJHegUH5tCprme0Y9i5QWE1SvbtfBVNyNrgPSRCw/J8QIYl
clxWtidC2fq/4WA7I/k8aY1WJT9cJ/GROixMbUvXJkMq8lXTm5UUg/vCVunUCWJNoxSRLjCqkfT8
ywDj+X73u3cAIdgm8r1yX4FK9ON6QB7njt9/2WdVVXVfndRgl9oQuChOmUr4KBAgsVl0kEch/A54
V/1M1cI+YGzFhtOMxOSP63H1d//od5Ktk4Czq9AalABIrHs4Uncz5N5+bVTEeERTGsPZv0ghkfkM
Wk+74jG5k0Z4K8cpSVaIlxauaAsi4eTTmDD2gIN8YCBm7m5fd1raaPZ1fLOf+mHy2CHmQBR7b7mO
Y4XfTw+wFLC0TVZnkWpt1/mvXAkKIO1+BNS6km4KiE54lYRUxiRpybVb67kz7C231NwA7fEHuNAr
h5hZtYagIOe+l8Hy8hmXf30VwHe5Wh9RbsH8x+Lkts5XhSSQp87CZ6MOEQDwFM1D0Pirq9dKsAh1
Uu+/xziJuYOIPCSISKsHiK56obkUdW00n1FKqO4HPQZ6Ki/6EvpefjmR+fNDr1w/BRcnNDnxq8ph
b8SktX6PxXB0HCQaSGJeT5TJCbsWHUIOsNxZM9st0LtDHvIMMRgd8ctetq7/9Mep92BrJCvyghQK
MfXLbPy5Tq+psOep+ZC7oPuY6R9B9ojBTeeXTqUtyik4n/ZOOy3wYqMh0jdvwXcvPGadhanAJrsx
gPig/dGd1VPYxLUb+ortxrH3KD3T/48mhbAI5tzIUBE582FR5hfKo1+7h4nji+f8yuS8RGXebZ35
kdPb3sxpznhFWoymyC78PasU5U4H83a3iKYe9cm9mIKPNHpknjk8yPYU1Zu6emWIlpIkHytpOwOJ
VHloXaU8e7HvbrF97PJdU3Vuyc8OkYmfa7fQsxyut4y+Uu7V5BVfuhsGsSvaibvKI441lYM0JSIW
eIylMXurPjdn0+TKDewfV/tBmIvw+huPaUOa/o8iOlxpDEsy6FOkVmLL75Vy2wLmon2z7Qi7znDE
7HruyxoZaC77eamKGXW3QnkxF6DDf/lMb92Gap8is6/JpMQYdS1B0pOZld6Rn0oEPxiaQhk/B8S3
yE04AfHjiHG7mavyrpuSwQ8j7NRBX3BFKvTfkU+cd3wEvoKy1LdJdOe+ltKDrq9uN3irmIvT2tRz
LAWV6tz+MISf4sqOez1sMp1LfdypfjSF+wZn/f/1f1zTs36DCzpV7Yb+vO2xrT8t0IieE/Av1dKK
C0YQktTLw5Zgl3M4LkVSfh2u3aPGL1Cnq2Pi8LB0nMnVCgNmq6WY9OjglaGI126iWKu05CLRpVkY
VP+hiSko2MTuHlYnKfysLWg+LqvEEFaRD55JmIM1gdEXywQJDzVGw4pJmlBk4rhTAHphBnRorC7T
83UPEYFS+fU/Mdh3iutl5HpjVZcTyhDLXhG2vbO8XTEakUoLRWcWzbuU+/BhwqFArJxn2ul0w/aa
Y/LVwEjTo4Fa00vqTUsJSz+ZEBPx9R9XrObf2PnU/gcMCqeJPKpck0gfnWUCqWSwF6dVimz4x7e8
fBLYHnmuw6Quz2R7gnluMdURkLKa8EnjKhV/Wx+IZHRZ99Vix5SOvrDziygx+F2YoOvocJEDjXwO
UxCp3wgaK8v6AJx4e40VaKDhN7LV56mRmF2b5AYqtRGxArNMOj0LN1W9xkkPo7e36XjrK1551vIy
EomepyLsH75E4hJxqjr74IFvkMofyBjdYJ3pvUvCNMPHgfrMFh0TL56OWtBl7XdnaBSJqfSBYRc6
AnJnwZNjC6Bd78Ebj8qdwnDNhTBXxrxuzTDlN7l0mbN033w8bPnP6wFYYVO0dmJOZPNdXUVP9dql
45LSC5apmgkSpp33wxDYk1dIFzHPLRt1uZVo1HPscNLxru+oL0lwl9YUMeXR/2IQmw8GcycvlNYE
WVwrD3YobGgdpIISs4H8Od5Dba8f3AuESSzQPoFZoJRAugq7j7tWHHZcsZ+HqWb3iCyBBR/UQB7U
Wzm8Vc7l+l/LpEx9M5mo3+h2/+ZhDmJOPr4hguP36moxA2TJYn83YuQKAg36CVMVV4tGOJk/vpt/
HXkBSW6EFtig7I6AsyIE5ZbjnSIrNtW8Z+HpG8qPyqQGgoBOTLQEivnry3b2Y3ir6yR3jF2/Y8uK
xeFy3QLPbBOZvcJ9beOvdu4qbqItf9ELOXH4j+zm9skpKARQ3ppzpnIEsX6X6qQJ6UrspHvybNXf
lg/y0wFO5aWPZQIHUoWEyYjY7A4Va7q7h6FuEqwl1Vg5SDCGv1FdPeFK8Ddh8MWXg/c/uANHkzPL
WFRAqYdSDQhbvYSVvaENLOOsDBfaXHP0CzwzC2wz2UoIfeM1rtnLJhTB4BI2Rfs/JiZ32gNUeJ59
LxaDu+LVC4FmvUY88ogfDMOaSMGkbkguyeaMQIJhzUgPs4BFywR79Q6HkuwEcNunKkLhSgYYTflg
4jA0w7AfhHEVGf56uum7w6wIyp8NhdxV0s6sFZwKDqu6XXDKFJv5xHNVBGI0WanWbjz0cmMgAlBU
LX44pjPid5uYrz9pVdfa82TGbHvKDL9/bjfjpJSqOjl6vRRsdgFSY4pXzoHNsziirLZnhDL+6YdJ
wNMV0cHk6RXzqAJ/MG3PB5nhbvlxX1K71AsJyIzcZ0snqpQJ/K8PxjYqR3WjDsU3FTEseOQjg2N4
99Erw5kPZwAhDsQ4hgkac23YX0//2mIh0wfdXmpSTW+atW9cKqzkVR4YkMzDihjOMGcq0Ikulhtw
hxk8V8RJugoK6uh3XLRMlyqwrw6ilkewzKCeUWtRG0JKlP/R+JrDVQ00pXFNn7FIJcs2bUCE/iV+
nuCwawpgg46EnbJsQYMnb49vBLluqVtknaBjHUEGtru+XwNGwnRF6LiwjwpZGNoBSJbEVmrfsWu9
s965isSPeJD5hVtGl7Swb195iSQoI7y2n9GnbgQRtVCZNAAWZrqWLtMHlRPEkYorIkWiQCnyZvW/
yG5KtKqsOGgI/GCHF1gWfYgWKsyjPSGwcD0YYpWVd/W/OJqKR+jNFbJQpRrC75vcXrteAO4byQnI
+siHiss2T7WYR9me5wclWOTAXtPoSNVd5rODjX+2A2w7uMALXsgV2ntIfPyFXMnJrN9hQzHHv/Dh
JYRfQ8MkVQoR4bd/rD1JvN4vH0V7drbKBIrTm29X5eRFnKYWeVLCCNpckZlDFJwa0zDTMp3Uf5sl
LKT0Z2Bcum/P+qJqqrfbE/jXQuK3/La15QC/jYgCDGAEmNm+7XeMcpF9AI52yg63EMb15Smes8t7
3qNEvOpOKSyh403j5j1Dr+soNPiHze/iYiENc+nEyRM/QkC7WrM5+MtPlhH3GHlo+8ETrwaKOjdF
blTw2SLZj6tzc8SQzdZBxvt1SgeM/JUwo50+PPlpOEHgMGu+apEDQDn5PG0uR8QacMYQ5lRXfO0l
To3ww4hcndZFSvuSMklqmYQf+pi0tRkpC6ki3A7Tvq+92A5GNtoNXg1RZaX9qQ+VFgw1XCdHYQs5
hxankaDZUMqzYmFdWMNf2n4TegllLCXM0UI+xiDk35fsSQjXD2cDfqFZzMnCIdZvHBDX3vlvG7Rm
nKWlkH5Z/CtGi+axVqN8dFC78Sn/ZgKnufyDfAeF5j4UnEv7sWe1r4b3EM8auWKy+1OCV2ejUaGD
wGKTCVwfH2nWjTBBXmX6jVDkjvowD057+FKsZdYOJqfKeb8nof7y7xyoUJxQ3xwA579cb3J7vZCq
7LoZgpGuZ9Uo52+iWxOQVldnCyGWs4yaNFzfVU4iXBDIppse33XFONF1tANjx9eo4iWHJQOiMK4s
sZNayZ2pdN02BJquX9CjaQ5fh/2rKfBStZTFVrs8gnknm31r1hXxy2ir754f/KrptV+EzY8uQsp7
1eTHMbH+jDqMgLLGv+bmlpCIhLhaxn3oH8oRSlr2Hm5mDXHeN+pCZEMmlNoVXcK6UJkZhPlz0UZP
tHGtDr9Q0lkisJAw2dmGDJ7qSMHmZx5cPOau5kNPKDSTzCnkSdhQ8jnjhm6fZIgPs13CUr+RwYyt
MEh9wnnH9Bqs2vd5O9T7XuCSyYjvMAs89DUvvXWm2P2JiIDKfqLXONMASF+fm008Ah7cV5zmUaBO
aMPB7rUy+vZMkze3e8b3bQWgQDQ3cX0dAWVxbtiMwPGnUXBxu6NnRF1Uqh2EE9Wkq3dHM0qd/xNN
4Qr+30mjOIIyaGsJ8nXOHBXVySxlU5+LZljq4bgmeVC0u8y38K/EHJkrWnQy7SW6xoX0DsC+pe5u
uK/ViEHYyDr8YoFL4hWUYKfSe3Y/yedA9FSA0yWmFoNYH2rKtTgZeSi1L5Vd40u9nn8vpp+5/H71
GdHl/Rm2BdDgg2G7KMm6AT8Yjs0e1VgxtvB8BtzcjyY47BnmKyamBwYMG4YpgexbRZ2r6u2VqoRd
3ThRwZ+U26TwVDXcCLi0b6WX6Dct1TomYtUPMUlGb8gTxC+OyBcm1w6aTJPSdiNoacsjGBH1/EZr
CfeezbtGNhXT81i0hDXDVwzkWfceCtFdusW5DeHlzbkcYaU1C9VGU01j5rwd/p8AdL8W068rXtm4
WwyG6HNN8Ht5qZ1iNcJqKXFjGsnRopHZ21CnJKtPsYP79TktXosbzpf+WfP4hFRQwJ29TtKO3AVR
lcV7VYV4n7qHRKgsnqChlMsB3e6+clulYlRTsIsqyNcxyMzolziIKtltA0lsrJLH4b9Ma14ftfCv
XFF//Fv7GMXBizkjPyma2ndxVEM83oxXmZyvfKNJ98m9OzGaIehis/ex8JXsXFI6VdcByEz6MKi4
yk0xfahOrFXW01DMe1moHRBPW4UZKed1JQFMu/7QjeaM0MQ772WfIfY+EqwLpzEpUSwc7pWhZtIn
a2UL+Eybj8QgbgenGi4y4NelcsqhJR3CAnekV8gNcIuEnEznb4LckFYRDqlHPrdz43L4LU0UbZyE
xlYt5WYHwoNqsyAPjzwCoKWVPJMXc9ehXzxTLs1bX+cYXsbNYMWKZqYmgt5pGAEatQ5xDXJI3Fu+
7xwa1F0emlvBAGvQw4J81FWfZ4S+9UHmP13POgFUwo0VSM6nl7hNsxS039j4qPIT3cly6SEr0fs0
JlalR97UQSJRwZ4SS5UHyGLSgZkE+/qNRyYqkOUULKCdK2GD4mMWDdxxqhhZA0gxgRQjA4jimU2l
dyo9DRbUF5hvXNvZYoAS9b83ac7z5OVJ8stI9+l7gaYPYiUkBTNA07M/d09JatzBEiQI3DaZZoMU
IT7JeA0wXGI8IbLmj/5cZDCq8IoMC6C41oGmW2I+mmuy5L38dut1AqFV9E8CYnh3xNs3hKU1AIx2
9WYMG1Yl34cb4K0pGzsm9C840adMB7sM5normAQotNxjY6TMaY+FdZ1hvwiIUHWlU3lwvneYfDpf
VSHPxllNFyhiacJalqJB9PE6l/9Xu2Fv0INAHdyXFKBC0XXRTPNX2vN+FH2cpbVa9EFYkTwypAzq
mcHy3NYqp7ZTvB/AEh7DUxRcNq4NTMVmJ+1eVnCBLOAlvWOkA+6FiObfdatO7GENKkS51KPxG9R1
PUdWwnEoTTHFfwK7mDHWLegMIlziteJvjykoOPbD10XKidkyypa2fKcKVr090UfQYwH8+vk+D7ke
dzGt++YSHC+maTyXxyngnc7G0W71L36U5NPeDUkWexTP0Yu0uGMX9CSAKFRb2a4vjgg494FxAv4J
hPvo+vCZQYcNCHMuofzZGFczaOrBP9RykIN/ItAAqdOoKqlskl3S3sbNVt+k39YE0IuV/7Z2bwc6
AieJLD8KiH9SY2pMMRR89kolUcu0LaRWmwO37Kr+FNDVYYf2mOSvZL58YCCT+w7CrGp9SEJ9B8/q
Cjgx08ycld2e2THs6DvLOmT1I4IxRdLizcmLj7M4fDHbVo5b1dmALgN2rRReBhM/fG63dnTTms3D
RT0C57wJZk7xHhrL+tHq64Wu0DnP8t1khcAeARo/+4IPCBnChAfu4p0kEzn6jXuBo+qr54I7WdP3
6HjaE4MaFFJnuuQNweedql/B0TEzRNRvk92mOfOhCiI4p2slliaApW11cyszcVUgf7+LQ9lWk0/G
lhPGmK2N/dJXbvqpK4manwEstwueaFTc6xeSbrEjBmpQAdAC5FOCWIKvv5Z03ecJbNFY30I2E+58
YwTEDkvMyQDOnseX3VqZFXxP5lvanIkiT4iunEpVtSz0DGBuY3+NnbnGFaIUdXVrAqRr/Sw3vGX0
YKl8E4EweuWxb0zDiLWlqEZV4/WlfX7a1aYN1JI+Ly/jHSthYgU6Jfb7dSV25ZvNLdYvYQzYbGUC
H9OOFAGCHIxfAIfBEUYoKYBhk2xPgjdb/JeNYUEQjKIn9D0MGxa2RW67F0rBxc4WG44EhDXq1y24
aIDvXkTDQ6JLn6Cwuaj9PcSx4OKtNFGJOaDny/xFzG/i6jhLRz+om8c0M6SoL+XZluYMaWLB7Lio
1Cf/1HcpePHPak+SwyBMt/2aP4gWf3agK7W8nDQUQMsAhxEgvtNuzxoo98bS61NL+d3FLHsoi5wc
OMIu235QUfcIc/o3VDYvezPcLLl9j43xe/UxAuMnAWNj8Hs2KDU9ZC7yBq/W0YHVuS9vELrtFXX4
0M7c1OgatiFgmITPaA30w/DtmNnHuZyx3DoXg8J1LyNYEmrLsdd2CqjftmZ/lY+uxnLIEQ3TeE3u
cNm2gEFjbjZ6EWFYdI0OVqxlDIiJIOZe/+XMO/SaZ/KHp2GTo1JoPx8IOwKkbV/F+swpTaLsthbL
mrJCIhHgBMxuSG3rRJAp+LZg34hLJY3Tu5ormGmWPl2pDvNMybrt/49DMpiqdGPe95UzjYVNb93/
kg+/LU/IAiTW8ecVscVsAJF2MpQVMRGQCA2DARsu/w9UxY9ei8xGZ7Rbyaw9VvzEDfc2bGASfcFl
D2YyDPXlTPCs0r38D5HFRIdU0X1r8mmaVoLbZv9aI/RR87TxJs+hc5z3mSVTMZju6roQz77fbHOK
lb1p3tZk86pKfuWOLupXX4DR+N1Tr0CVPzc+IdFOapnnCRbqN2e+zJU10N700+lNCrxZw/Iy8Zyh
/MiTL+OJ8Z8vt0PY5RW88cXumVu101gs8laQABshs4MkOyyTn5aibOqzOXKt8ZM6KMHE0+4+0GwQ
Kejb09gU5RCEn17jH5xQX8nsT1hyzoZy/VXhXZge7wmmdSlKigzqOEyktoDo/R67OlZEVt3zATNx
GfjyD5qzsuXfPUPQw2h9hwGv1mR3sVuy4XafV6bRYyZ5unMEVwL//6xOlBD+2sMpky2yPjl7n2pu
+cMw9SWTKKeWWGytUxphwNtIPktiDyypip8b4L7vFF1HKdYVtZ7wwy0WqqEYdCLpDBQ+4yy3pej4
i/4/0jlKjHb00sKIcwoZvvUA9Bg+1qbBW+H4rbsB43+O7OBpkiFWjMCJUPWRKW8AdPrhIiwD6WVf
FasUfrCEMsK/ayPZGxA19+0c0wuaQ7X79DpAchFPf5a+9cYyuD3zfiQ6wL6CKDrGLzaEVx2BXMEb
kRW9oeqfI0yo1i2L/On2cpxGL1byqokuakPBOQZKH+ASYiF/4q1169PLKtgrylZ6EA44ox2MS11b
o3w7B5YsGmBolW3TBCQgJkfJXACuEtkyzFiqWgcYWUvVmbPubm+9Es0R3FkzH1uTt5Jd/PJubUSp
zrE/LXHwdrzPqi/md5UIVyXKdGlAi8M5D+U11M4fFCjTDkx5kFR6wZ4O/RbWJ8r2Yd0qHLTWJ4V5
R8c9Xfe2cgU7pYmRnTRBfTKWuvVoV+nWzc1z5Jy/qRLuc9P7DpDLGhFTje4tli+iM6EAo6r/6/Bw
5RRdD4eaca/YdGwki/B6DzAsuJkLDmMB9kDsr2oOEki5Qouk5zidT12PKRO+9UcQap7/Ej/LZx2u
HccjrXLbtQs0D6jPWDvA0ch7orGJ2PxwjpKMH4MNC++xShZ6BDG/7uZCJcqbCky4d9XHy7xg5yBu
zIkNgAr4Ge0ap6ezY9WxSY/fPeYpCftzk3YFt9sChr6Mzg1hGLY5MLNsRexPsZdRmQ8ikyBIgGPP
wxDSjUM0YLr7Rx7klWvpDtS6EvSRlfMDlUS/WynLdgxSkJvR+GMlgSUXCiYxtzgSIa5gCrAckPaG
n633SGWU+DVl3wpCeKsV0slHGvNJ/rVZHFdEsR5H1gCf//BYV/IMVVhm0piYGMFFEGXT2f77wilw
PUso/jbkj4i9hh79HBFZrLiK2Rxmc+b31kLhC9FwjcERscgVuIdTnK8SaV9nbzOdKiQJN30bIxLP
raeBUzyeDH4b2lrJcPiO1AcN+diG7j+CD3Cy04YCK1rnohybJpjQc02ObP0ebyu4Ntfz/CE8Pcva
6SfirdP5rydAjC+w6Exbq1xadz1BawCcN6z3FmLtd9Yo43mbmtd2+TNzIDtPNE2fFvr+e/ODOfTs
vfu4StaoPnWOLWryBHG6weQNdwOrMUKf40OuslNBj90fQVE8t9eEwbpC2WYpKW9zM3gdyHMzZ5iB
o7QFXaCeqNf1Bgii5RODHomYXcN1FaHe8aiiDEAk6iXZYs4k2UiYdc2+Mw2zY9QhBSlczqqX0UFS
U4Ug/BXKcUEN+ft1jHszZHvllekKptvGUuDhhwpJDxq2XhEIhO7d4kTF1RyqFDnWwBwLU9MEJl1C
cDlwgnlbfM6Rq9/tj8yxXN6p0s8jtiU5fnnHlktekAwymBNO1F2e5GEoxdsbt67ZOn48Y+yNZOc1
qKVPpsypIN3noflr83YOVmy79llJo3MaZdKjcVJjrLV8RzXoIJk1aaOuO06BPZyXRbaqXTSVWM9J
reDSIdhIS+6fSz5zVBDMT10ctvaPacXiWq+l/Ck9Cqtwf1LeaD1FknD3gNoEUp6okA8LbuFnTJpI
N6zql3MaLBUTlnC4jpR09xKvJve9GDaURUC8T/PiwGt53a6ak9XB9Sov4Gfv68MsoMcd6zy9PFUs
sfMgQEb4iXxVDd0hcRVvukIDYGCmo9o8Vzvyjl0D0+YJ/UGbRn7038NyCcOQJNNlyMED0Uo0v9W+
bmmcYHlBTLejR+gHH7XU3NbY5aDA/hvT+VYY8Ua8U1GDoHfYH0EFalLyMhJQgTSieV3hfT/H3t1M
2v/03HuEZDkpJxS2R6I8lo+pqd1QMMyI7xjvGrifpkW1SgXzIervoKeXVSHUKEC97LR2SAW+Gg1a
hGNTyLWTGr4DdA7Zaw+K/bVKNDudswEgJ7ReaUxHL5mn05KKmo4Zw5x5IEE5lT7fZ4CL5Ch+6e5O
FBfTLKMd6h9J8Jd4IojJ7D9bTCrORtM1038+N997jErFTCU//Lp3dGLGb8XLK91QKJbijlDV1wjk
HanlpRBTwh8Dz2iVL0ffZqWetiLeMRxd1BN2/sf25qFoMMTocfd+w82wRDpfgtSgr57TFiTuPmpa
qsRgKvpnM+ohITwGRAhQ7jSqof3Z7uCpHXBT+LWZgsF3hcj9ZJRHMr98EWA0OYbZYrTi81/wgM7/
CviJVkLEm75WGMHnroyFPq0NzrlAc0OuuUwFBCPeehw3yFKrZlsQq4lzaH12xu/oEY/InyRO+Wc3
0kpHxlVLqwj9Xhytru6YSNrIhUgmWRW2CHBoZJwwEnWF04luvNIBPKi/ebh0GQzwrOD4wsazDcRk
e7eL5yhpKt7++XbIhsz3YfnBNHYyqLg+ivZFmOZcXautobIglPaw7AcPg4lneVK5DlrrdANuRnV+
wQdev9OZU0pFkIriN/kFGMRll9R91GHZmJTyC3r88P59ecmDhSHzItYvb6jEJUlfoJPRvsyLlnQz
X5t1jD8T0X5kImSiF4oUljXG/BwHtw2EHRji0nX+MoX/YuXFZ5MDn+uAI11JU6tOi6AQpr7bNnp3
SV6wmaPmVU9cHKAfv+jqHmpWjA2x5rxZT8CeQvezS/3TzR0JrbYI+YO2hsCYXUqr5M1G4g1UAJky
WYXjjPPPVyWnfjy9mr9nVr6zutZDygxgLMUDrV7WNNEHeTQFuGCIq5ySXgToBqt1K2duyBQrS04B
jAA5zk2o2Y2Akr6dtkTPtlPg0OeQWuYhw5VErtmYxcT2rEBsfH9WdpQ/QdvUFrLcjfex10LsIi+Y
vD7tzaExzy2XsrS8yLb+2dcgsdYHDTj7XI3pIiY3/DF2W2IEbQQzJJUp/oykSzD1sXNH3LNDwud5
ObP/uFyGvx8UGxf9+98RP6VtWFNLDI6N7leP+uBueJ7uvkNFRx7adD19HgKFhmnpkZSQoUbdThQX
YhJh9iElzWLorqkrLY+tr8iOPjaTRG2ihJgLVVt1yd8NccpVdjSh+SbiLS9D5MUlSVF3D2wlFiLj
j11/pa2Xu5PHLBLXwZO9O4ZrbFObesL0iJDZTdlVL7ZTnCuY7NC1D4uPEdLGYEjkbCf/ued5PTUD
FLy8va8CSCF+CiVFTLE7wOKeG4zZVJUYUyVFlitsRkIMr2iM1TqE6t/uG83oc4Y9hLoxswa72Pss
DfhtzHVQpW9GX7yrQZe1XG8bRZoEorfof+4SlKFsNCcdm9/UZX5dVk+rdGVR66SzIVoNWntzDIoX
G05arAwELAzMdFFeiIqZZ1eCL0rFrfbwB78c9KJGbaXXStEflh6XVRJ5pHo5peUBC8ytrPVp5XvT
g+4zFY1ubS7pLqurXYIUMqVo9+9ESvKjAg+ZKSIvkR8oj0DVkUA9HtQrQYudnt2528WFl4NFAcgL
TjnhEWfEe18cPeqC/8fOOQzSZLD3riLSYBxz/f7Ny64GC81TNjDmMLyLDQ8IZAQ5Amde6xvmeiXq
rgF0G/BOPns/kHBBMixYLXXclvQBeZt2mmxKhlFk4D8kujemHld1nU4xL4p1lAYn2yjPE2O4Vro5
pS6FrMhIkSqFo5mtlMQVIJ5k2NhJrSZT7y+ZBdxw3IYjK3Z5fPX7buh/kru56joz1D/G4GCF1oae
b7ztGsprR3+6G9tzEvvtvGyViYQHUhqOHyrCgURca4Evr74YZD7qaez1zEIVfwlp32P4ORSvOsUj
Z6DkLwDtrwuUSyrFuWNscT0Pa124uX/rB14MHpV0pUWBdWyONkpwlJx10dl+DGlA0wEe3Ig5I1U1
Seve+3oBRikUm2PgI1lnbYQYWESCEnGuCS10brO2rmLVI7jRcAv19IKyZIGUPFkUxSpOG9Pj+KKI
4i6QGYdLp8VSoRfHRC6MXhkBTtHH2hlXIz1CzqnHeMkKb10nAFAdaQu0ti655NgfVnaB/UZs0F1E
FzUXN+GRqvaxmvSQy+vl4DikEFUQ9FnN3im1LD7t0+17nUWhT+J/YGU5Vb1g41N8V0tGG+jrSJLe
dKCkA4r1CFXJw+05GLJFX1UOig8z43MT/9ZxVnApy+VQil7XtCZRerFNGQnI3h1GaNiLeXL9YS6W
hrjWmZ62w+lZRGLz1F8CzmalaPJfCdcjDfbEa48tL227xOG4hFt5YQjhjZomAxn6WotvgWHRE1GA
RnX+1ZwrjlQXoN52fAB+JKUV75u2bx64AHI4J59WENo/Fvd3eM2c5fD7Rca7hErtRRflFZtArnaL
IZ1QTaBJiKHuHkMVIkd0wlDOAEImQHbkdlf5ja/DI3k0ajKci34DKOddlvLCCoPRM07QmuL3omr7
6cdVfjFzmFvItUkH1e5rBnoGyXcc0fFC1vRsa3srxPRF9DT3k3kxcWot2wEBoO7oPKFJ6FSovDGb
pqcz9hztQ9tO3RzXAxDY5v/s9HVsP2Ivn8wzoPMyc7SLviaPaPmTOgQ9o/fZOECsZ3ZPSEuX15nw
s7XFYpf4LYFAWGmSgwCR0q8sS8BS8K9rxDQqTGE50DZYs6uOeln4JmnT07KwjQfEw8tQw89IOZ+5
25D+AhheVyZQSZPw2rHRR2Fi7uQ0SrHIHlg2JPhKJwizoSEN65YA8VKi9pT7K7+xB9tQdOdDcXNm
rRT2d6IrKwB5r8eUNhfsPskkok7OVe6muuj00NSDQaHUEMCR4d2DbvOyPLnctmcaEP8St5xKrJyk
wZgxttm8m8NjcFYZOaaVLEGaOs3MyXl6n6HAlQmHUpU2MpHlhOwlsJlGQRYbJVCAK6kM0XekevXA
goXMEHG6QckzJOqHw2FWlqMTUvukt3QT8H1QP0LAFknzBwuZw+AIcrXgyF5leChHn5BjB4DTH/Q3
wnGyFfwCzOCQU6m4CosJgJZt1cIW0FtVrNkh4PMEzsznyMvVFt0Fv/wMMznpyjplatkagzXvv95k
xVfHdfIxFYjuLJqseg2x57k4F7KsP6GQAL38Ftq4aCFBvYCp7pzkkO5cO4/j3oW9o4v0HQWDVlLm
KRn+agg0nZdCSmv6y2Dawdy0A9FdTVFy+nVwWNjE4FmTXGuULTqq8cYrJ1Drzy60MgMz5hEaXyDC
pNq4KR8Kn3imzT7fgIxsuKemNB/hx/4sd664mhgUB78Rpb/vCRECULW1yczKGYbZP95/YRBvc4E/
7W/mLsEQgqA+Jb3Fq8djpD2g5iOmCzBHrtIQh5baol2a1cfTZXWzcYzOz1vCBLRrTK/Isj2Z+Vfo
hyfBLT9DXLzFLFFvelSoxMfdqSZhuFFfQawiM121+k33yu9LT3cJWiFphyfftS5r7Fk9WT91f70U
H7kFT3IK8zBdsqYLgchOjB2DuFXnjdaPFAKPld2xQPNo+k+JUtw0yuoA/vXiU2t0qflN4apDtNHH
sA+vrwA5CUa3HjUOrKlywRSB2IpEJfKr+ecctmD85KZALBD2CUV+c9f2ZfCj+IquOiZM7PC5jDhq
PcMdYbo4upEfpEmcic1y0h6iWBsKX6f3gZcsfdFAzUNlG+cQRi4gEKiR4CMoruPZ+T958zw3B6Cw
DwagsyvSGB4vWAqT5HPVvgVaFAqoiTPr8KSXk9FqBDxh1HBaFAnCquu8vunnDaTJH8x8KD/iPU93
QvB/ICqBmtk68/EFa5Bjvf6+vxZMn7UOv0IMwYIAuMM7Ws01dWeriKztXwH4pBtUMedrv/ps0/tU
1rXpewcgLvp1Qn8mlZKOeEAln2aKdUTmgXFcdU4KF+ivdzFtAXr7u4idju/CE4VzJuubYkCNPLfn
1p0xfkJ5nevLrd4mF0V6mzCl4FITXR/KePBIH7epRBci9RmkBCabC6MVJ2JWCFFF8Da3s5ihBv//
jTb/bq1iEDHiyiY3tdGu7FS2Djp3XqZCNhyhq5JZASZQDHa1aLfYT/y/KHahWCG4ysL0CS0Zl4wP
JC/+4sJ5rH5nurQLpyImifxs7HKvhJcP9vGgzmj304ym+6KN5RCPz1SGXoSm+V9oeEcfi1KtovCW
ZckWK9FJxA+NtPEcEvICa2sUm6Pi+ouRX+VHpRhHRci3h1hqUDVfjIxVFSBUWuOsIzjQ2CbzAZaF
sORFvO/64N9opHcUg33oWeVqqHM53++5h7kTJZJFZd9H/npgqAP0OfpouezBU/liHHYAHodQcWRz
tI4gtqbQ0J79HP4NkuV4+JyFRu6nU0DGG1vE7fLlmMuhgDOVDl/sgml3i72k5PA/8aSMuIy0P6jn
7KRWfPKQGj96LPQhfz9x7o6HXScTLPXeDTzG/cgFBpn1NZiZvdvw9egXZcY3iA5YhMJkGFCQeVar
jASUGsm7y3A9wuJ3oO7jDh9E6jk6vg4I9aUFJ2bImCg224v/LSOTI/xEbGml3xKpkiyEQQ7HZ0+q
VrZ45NvQlnMUz5UW+MnTuHl7qQ8onD7hf+O5M8dtlzt0sbdz0wynu+Uv0duyo2fjUF9vJNRvBZwz
36MGODWRuDISnp5Aq8RUXhVAh/VAYPWcTZLmzda1DGZDmrT258wM51FNCqoLTeR5NulsGdDYlhQB
8s2Lx23P1oSKwXBHIyNhMNH9VZp8IWVPEay5o45x7kqzsuUVVkNIeCowx5s2am53yQ1CPsYWBQTm
GZPSh7WBPUkUSdTbRbmGc1wIy+k674W+3AjvYQ1Vy+mTAvAlKHHkaAMEfCjE3rXZwSYTDvErpD32
y0lVSVys5xSHP1AHJO7mIf5mL1GKJT57Ix1Y5drpEaztQI7WSXhfB/I7CnZuNybOZA4SCU3BPaJ7
yKyJLTIQ5HBiiyMe5IfqouchSqHjF+pNSG/NwTq04jem1vTsjNHn0MdG2BdcfVJHGKSCJbaPT0iM
6GnvMihw5BK9bktCe+Cuvouz1D2pHjNMoV1OEjPsvHqr+FtYD0cFk/p8DRmDWoupHEQQADxtcLXS
eI3Z/hgj14HPR5vU5WLj98nXyy7IHuQLmRLsBilaAiQ3U2p8t8PCAoa1Gm9v/n+9UkNrpN/4YRyC
gfy3wICed7T+aN7SsBbScgsPh6wO78/c0akD7S+YxgTWRV6eyKyNkHIiy+8divL6EI3/18SIUIW/
IuL5FPt2V1Q8PyA7qUDffKslw+tqe+nLiqfdE8mIcTmi1RYLAhtN5KiI36XmUpkMKM6u1L7wDGOt
FlVz57GnMS0mWPyX/VHBuxAsFuq4RnLbyzAi3KaSFZV8Lv9NsWtzZm206JP0bP7QEQ7LKkkaYbqr
53EWQ/lRTqeC3fRzafTXHxFdbnyxKdZn568oz5rebiPZn66pldaDY5mlzmTOlFDJaUg7MEjivfFv
LKI1TFrIwRyNI42oGSdE6v0sJSiK+3xNF39B7jIC8EjxK7mYXwJJfMNMBj4ydc2MW2FOcyBbh3K1
TgzeJtiVAC8Q8WYpozcJPCWcq71uR9+3uZzSLXUwyJlrB4SAGoOzGIRVQWlxHV4Qdyjud/j4dkEI
XccnJHjgDLbn3rlU0edf6oTTX7FgfbghmPCcyD9r4qQbMohNpISEDniGpNadbf06HQNas5HikVU4
VNMi4OYT8j4hHx/fM69i5hYE5nzcvKfvy6uySBdndgPgE6Srsell7sXIs6bN3NObUGBxuvbgBQTl
a/p5FcD6NDF0OG4ZpkWyI+RFcVl2uadn2fzMRlqFMzu546El28rdRqxiEXc5sUxHASth+Eckd6lX
irSy7v2BLgP68yoJp9ypzJ6/wtNAfocLiRCBEGQxYYfeDeSk7GViHoTkrodfRg163hzy1gW0VEd1
fPColOzYMdHtZHjYGynpBKMXYrzfP+ibrVnhZ6CvOKXyBjygPti9P9LPzLH6iyEb0isL61pEqLSt
WgsibiKK4P4h7DbYrJBDbLc13GkfgPXlL9fL1F30M+xZwNw5TU3l3jJxhZDEzyDSnxkg1QUjD5Bk
Eh+9YZdxWfxJq5aHrIypAPjObdg8S5SJLa9GbFNoxrV9oSLF3apvnskxUK1KjjpCxUs4++6KeeF7
ls3geJ8qJeOw2X+31bWi+9E3Vi0aXjDaGjpyccdpGifofOZ+LbZ6zr/PtTqKMsfSP7r3NbtGKIXJ
4NvWjmf2jQaCNFmyBkRfpATqC9UXOh4hFOTgoNasHR/0639DTaiCWfVXAwQO/SXscx92vqOwVVip
pKcX2+55P5QXOWFuOvpJBznxAWbDZMyyNOTDqrUVsvXu8zWNTOslOmmWKSx6T8Ac8x9XM9XtwlA7
uVH3WmHqskCUo6sezACoqsw7E/efq3jL6PQWunurnXOAwyZNWzF2yoS3WKQJRwyqiiHlzM1dFKOz
8t8uAdK/By7tSF/MAbbV7ST9M3/lEcuqs+EkeO8wkL7M60PlMHfnqDQaoQGLN8zN93bzynOysVxx
5uhG2HIJ6GHp/VQep349T5BXYB/G/led7Bq5eellhZTezC6MqCyj8LfoZ6y4mVBKPCnbbC34i/Ft
sMG5zGyc7jCow+o/yevksCQ9QMiZZ7VpzUHcAGVz4ZyxHWD5EzyTTTV4WVwtwomR/KWtGmL9nCFU
tLNp6ecjGIWHEmDOvITMyD9h/VIoY/2PiF3LCtlwNF4HHaRNIaKT5GBRZpp2BXzWCE73BdY17l1t
G9GImzRpKn9CMShwTk8O85wUih3bpb0pIz9Q6EIZzfTLEOSFgxYnWemeI2GCEQ73DR/jx9+QXANz
ijTu9/Qj4haTJN+wdv1YWm9kY3Dskdg09PwNFEF9Y4UdqKPDqBKwjPjP+RBgyHKz6UTmIY95CP/T
R37NeHket7tDWv9tYOdELcaIOWXrBgmiLXOgslcS+rQkP6fo/MW9gaQLIfRjp5Lr8B9MvqLB2zzc
IiFLxS+jQh0gl+p3/zIyYkyhTaMD8rSRZK3gLEYpLhk5CdCNbVmquBu/lfVG+2t5DgebZaHy2eQU
kGuUSzVq62DgKyqdzKOP4iIlKHQRJEG1P4uOis1EOQ6oIivX4UxqCJqb4NtUu3ap1s6T+JcYcrOQ
qY1Wro5tAdJq8k8mUagk9E2OE7Nag43eSh4J/w8Vjagk83N3ne89cuVamHvwKbiMhVI1zu3CXDi2
bta+HKAwPGxw+38OMQGFnxfWrQES9d0iIG/moIK4mmU037VdTvME7nNaIHekg70puy9v3zFPBad9
CmNHZUeIACzBtVe2WziCv1jcMeo5JA5hYCoYnIyybc9uNPmWPY2ncKhyk5a3bmsdc0Y7G/dncLW8
aet5aVNVGp8wt2xNBoq9dd3cOHI7rpB5Tn065xKtcl9LeAkR7l5uka7pm7k1mgF8xrsZ3SJlUJHZ
zWvqnhlHdOGkodtkaTU0Ho58KDNBzQO1Ff9ryUpP7UXQZzOMOlu42adckU2jDFXk0DX9njwyFxYX
VUxtjjxcBaj29naPmmGJ3xWbUn2KZynPFKDswRPqxwgSv2LI/k62p0CR2uPoPNfqFUCNU8EiO58q
X7cpEzwCBTykBbC8aZm2+4LCpsgUZhGHh4Kl0GrY53YLDrlNJCS1WSkihA5Ljl8eDFGXqc4FU0fz
qNciTXrKM2YCZCZLexjrRRlfp/5wo+gS2MunntEZIOlbkgMZp2cvqVqWZDWnJWVUisayLSWA3hs6
smPowLiRwOIEud3Sfp1Ep5wKQtfqp8HPXDF/J0yH7zW1eFgodxpRfx9tOiXI9wc/DIF04yRnVVIa
D2T4l3nlpfqwEMy2UBAYIGZBWs3SLY8uJp2Y9BrKp1DguMRCvWqsrTICp9GXmsiLPM9m8iHDgCMX
9elWaBU4SgZFNCjD8mH0N9SjXHLkVRElWlEm3XsS/6PomVp/ysqrQkHvOF3fotz8ZaJIT7e/UBE1
lSE8Hvu+ddmpjLfKRPomx2BnHst8ou3O0Q6Z7OYthVaB17xAUsDBjn49arCoa+9EwlsgColLzjNR
zTWmrKhzoqEFKspCUfNdGxvDRn4OoP6nzLFXjnQj6wFUAkqftqJjUv15Ikt+1H/mKyeGtgL+wL9s
bFNLWncgsoRP4B0839V7AW5Q/Y1tjBjJLJbnNnKkp5/AxRGIWCOqvN+LTLG8RDiMCPYqen2Q3wQv
XeaTHTb4LFK+5uUW+xXIRdx/aIxjE2qQYTQI3e+g/uSmWiLXzD0xn+7m9ZY5r4c8LVR6W13Sx01E
sNYBnL1xRxvU1M2UxD9yDftg24F6TwtFNd+uu6yEm0oUh2gdw8n/KAPPGlVyiFdT/nVinnn2Bsrc
DpDfV5FByt479/OohVcSkt5GmQtbGSIe7oiNDtBYuZDVwTKrFcWCqCqVYOthULarSheEhFnuDaO/
xhc97y5lZVDDtfkWq2/FAEAlj4RijVqPq8ejEVs8ow+R0ziZ/saYPjjE1/ozcCeZKVPsNz0+2JYm
VFii8pKlVjb+xhl0nctAbKEQ715y28GdCi0RJLQlsRS3s3lYivOmWuIM9jWOurYcnhsAfn5+lAJE
3SeJhMGC+Lj2eOODIUrSJTGWZ6T25XqlNJ3c5AMmYCElMXr1Tv3ZarvMjQNHtFcsxci6CSy9lYe8
VdTbd/kKWoQA8+S75lRw3CglP3KyncQHmu+PdGjN0cgPMKFd2N7aFpYwOaNXF78IcQkkySAvnonO
MZIhalS51H/j9MXGAoT4jeokLg9CUi2s+qCdUajttZub9bN1TEUJXHVf5MGfZYWygm9AFtpILOS1
CMEAkZ7NPNnK+IKX95mM8UNwFu1CZHPicDAuHJeVIQz44bfNqTgr3PhvkUrQaNGpCBKEf9Z4Ro27
SS8RYoojzn4tTWtRbSzKW8zlmemgd/BJcSaAlOlhmPxwVbwHEC2UHTXvYrLM0rNhfFiX0Ceoy2mB
I/DCtLx0h6kxeAS97BFh+HCtFNY4KgSZ+R+e3I2lR28y4wCMu1KZToCzoB9wAo2JGBrqaGCPihbG
rl9LUuqS4pNsDGQV6rsF+gltHB6/Px+E4kBwpsnqG2Zti6tlyyhqM64ghjVUoeIwczeL4AlpciN8
oxQhcMw1+CNV99TTfSZEdd9BYnFuorSI/2DAzFRCEqNwDO2626MVjMwatVS/on3n1dmIqtKKDC48
g+mct9YYBKXwdiCNq2CBDrC7QZPet78ZatkRDNG+42NLv1HT9OvqvSxGlfrVBW+zCjXh4zf5K+Jw
YwfqOEiG55hiBDyxuVzr5KoMZAgdhVoUzn1PzZLSmULbkxMI4/Nf611AgILFNBLC1u+DkL5Kkp+1
R0OrIJgiV5Auw2tYP4zRtz5N8cs2mfjzgMSgcKLeSqktXCBStG89z6g0g3g9r646YdG7IU2GBuwK
Eh/qJmDtEoxe8BzpgQFLdKmRRkKboB+CZykN3V93rot97hgFm3ykQxzsH7+KCCPHU8JyhG9q1uEu
7oLienreGX/4G6hume8edV10Ho8h8Mke0I3QP+geVbk4mzL+e5lr0F8iO779TVl8V/emyZ715PJS
pFWQMO0UNzSPlJAVi/rFj2QxBzEHCqESw2PbqAyPEfxZkbXqw2oqSg8nkmMvpIy9hfWWrsSh1ZoL
S04SBetOVpIvnswI6Fyg4xeOYFQ4yGP285Vl+R2yqtb1w8ENY4YEWNhf50dN+KsKwG8Qn6ElcguD
ZvFqT+328TEykh7OmPgaPoiSBqf6gIEW+EK4RM75fLvQI3tR4HYS4twsvN/IqRfOswO/8gz6M2lp
xZ0/U708uCfprRbahpvH5ANThdXVu5VIr9gxgYnTlroYlc95FuAgDhSTx/ARvwjv0zqpf7cJD+Tl
NSV4/e77no2Zxx0/p9JIvdfSRflgSNdX1MiUFFkwnzyBr1+wG6VfGTVxPSi68+GRZpH9n6G6OJS3
IZP33Z6et0z1j6KjLhMfwPBNiudoFk60dMV/PpdBRKLxZPAJlrra/tQE/ZRx9KwFYXaOqJIbit/1
RGLWOjdUm/BU533rCm5c5cD1Wr7k6BduhJNYvMkGNJB3gv3UOhagHPgZuI7aw/W15xWuORU8m0ZC
dZdmXzNxltzW0X6jEy/M3fAylzhYHVrXBRJ6eldNO7GdHx0Ud/cyMQ2/rrt1VPFLlsV8AWCDkl7m
7pNzyRhZ27sAuYR9Cu3ZnecxahOh8MtZYqdqxgniJOg6FFjoOhO1iFRVIBrOfXdqECoWiyzRzI72
9iG6CH270TNHi+lFOWYAg4hto9oLVdmXIikk2SbPfAvBu0Oouf2XeNU2D3aiI0HVpLlAtLsyRJEL
mrQ+D1zCKPluMoNp1x3BNc9N2neohN2vdh+P9X3zx/rw7s/26+oFm64RvCOczke+yZq4J+58MxOB
1VMu6fMwcRhFq9pnfvxbyRJyA7wbmT7cHYPPXleXv1oFwiyeFbBrqQ22Cvi8blCa0jGS9Ha3QNrQ
EGlMOfG9irkqab068MNLURyUry9My2WBY39EZC2THUhBisSU0X8KFLbpHnEWLUuKsFid/kUl0mmg
s8N3kD4+Vfujb6MYkFes//IF++xP3lHPp2P5iWpDgXkT/7W/7lFc5Qw9khqscShSEKIZ5FzH3Jcc
DYNzdpbKJgzZjaHUqitMmF6oazF2fKcsUPclfczuRbqT+Xy20wmT6/DcQtSwhoc4PmC5suYfcqLM
eID+BjeIssicdqVLgiFbrpR4xUTWYud8Oxf9JbhvCoEPE/ZCVZVFJ9GPlUqtNDxWS5C1RDJ/98iy
Npy5bTKBa4AR6UkzyDZBMHjftGaFivV+/DInm4IKrMbINPM3r1unSSJXQXJiEQYCncsd4HYXL1GT
fgxQ8bU/4/4crHeefNtsO2K8S9szhwpPmJngK0gQHvLh0P4NjXIKe32grycuCq8COvvT0wbWxiIZ
Z1texZ9BB3uO81sK5ugDOmsbrS51cIRY3J4FcPXZ6bEj26ihStTVkHoN9WKOHlO32Ldp92ckWXhu
h6t5AcKIZJBhOMwHw+PUNLqZSmhgAQsQ0CJIgQkXo6hV8S0KoCaEik/L0usG0bVJuS0GsoVAxHjx
Z4EPLdLP2zd37ThbpntDmPafSxOj5XaUn/U5WQ8kwKfUYt8mr0xr7TN3gio5IDXlvmf4257IJFjp
sIe9lrsxPf/npvxH9BkbvE9FSq1hYwFocpAsLzH71nSpia9+XOgd3vS431ivQuLER8sg2WSulvgh
fsDBJwExzDcdNvMnOLfYenVEEDW33XNCCHNjSi1GAOzKWjya+6a0hz0g0Ek55Uma+ScQVdWEON1s
ViT83c2OzclasYAGG8NuoYwZ/Qh01Iw92Lw9Tu/zP1pl1JvME33cofQFjWcEUyxysLT6/Y3XieRq
mm91TNqiGKTnrLTsQ4q+PFPVDbarFPlZPS7OFcufdEqzZgeSEZEmNfLunEn4y3S6O9OYmHHKYBZV
iIzpBciDbJfRuH6QuWg4DALt+uuq3XCA8f83GEMydluh7MYensGee9JxFHZZ1yn8VFGGVe4CgphE
7s3utghIt+XmuALVf3aebaMWN+5961n8Shqbr5PeiGzfRzodw4WvN66i/BwrjFYg5mK1g+q72ZtR
cPUQ99DLfSApcBOtgOBPO51navTUdlBGjwUkUM7zN4Eo3+0CpEyzTB3ll125xxSfwJPXnAnFuHun
PCx/JjXpIEQDwM0WdVKbfxeCS2TvW0lAzbAd1Z7Y1wwSkjo2MZZXn6GASCYu5rlttV77sIzyNE3V
ga05rg17H3vUXhnIRgheXOq5zEq6RAu5Wci+EeNxjRLwoyIHD79GG3jI4ZAdhhGtIc9QhLlue/uZ
bU3otCrF2juZLIYk1LZKLweq3fizqPaAXl8Rxj/cdqeb+ROOCpAzJ6U2fZzi91zTP1QPc9dybssX
4DQgSpF8JEh33RkR82AJQfsoRLbz725Snd4z+7LBX4bloFAoju9JInWC2teX/Rr8jVfqI+AboS2o
7d3X4/Ard8ZoQxzTwbfi8dmFvjkRK6PWwOt6JHVplb7u72gwmPIFLKpmcHnTLU1gmqnapcH2ejm5
qd2haqLruenE0Ww8rm9K1FhZSQJYLZ8AkUKgEjnbacS7rVFamXGcBHPFmC4E5/I8eSuyxOOCs3dB
3aBcDdDEm7ZtGgtk6Iz7f0Qhx+r9IDQWoPvpFCU30fCL9xbtWdQ0uo2U6VyQxqi85qgj3ixhJ2yf
6Z+DkNiQtEIDJ/hMgIBIrY3v3NGlawuvKEir8Fz7uTNyAR2Ho5NQwciA3njjHY9dxtW63QfnQw3V
3NoXx0nbj9eCNAeeG5jkTcvFtNlF677FkbSvcdQ/QH0szkfvh5uzDkdGEcNzYWJiHWHB/xDA1ghP
gjX/Mx+BNjedDDsVcwIP7OtonXsq2ac5Lwxx5Z/4tw492QFZE/YwwAM3SbXjo562/8dxvPgroE3T
HfQmO0S46O68YItHwbBR6zS8xcb3ZwbGgxwi7KPPukWAEcn2b3hSUhiG5FDElA2wAbW/B1LSauqt
JEPxMCT8PjVvGjtdWp9/SUhyZ/gxLJ3PzUNeZPvp0C81m6enI1zjj39pQYK1NpY42AFAkXTVUclT
Khpt5LNCX7fGrJVmI1v/92tszlVXcGN6wKgKqjWR/35mHhRgWvwYti1fxHpb503EIxcgpH7DEZcx
BR9KSTyPMLCkejxxyaxNT5FAJWs5nmUn1BPaYC2M+glYUN+ymlKIRrzvz1yEr5TdFTU+DJBvf7vx
qeVP3I69tzIw9ps3VjtxBnswjYaoog6O/+DJaJOTWydh0MkjrtHKHOHlnNsTHC9GtIRouWs+sS/C
G5FmJs+pj+2ofiWP7weW5KuHd6ZmpGJwdrTQogXvmsNZwyUYbp98GAQXXQLailMCukG8x6bku58r
YlIIl1CfwAAiBa0ivojfTzhSBqNfGQM3DuIr3vAJxSzz0PGJitgmE/W6CryYsiXxjSexDNgmq6zg
6p6I7bJM1tkzRBHZoQzCQuDFIiJdAlZfxY0Wm5mcJIQtEfU+Fhz/WDd6shOq5eNjJ+swMPG3GxAB
GTXzuv6pJ2HTlasV9it2zV/67b/Hc6Vh92M4Jm83j6tD0bFxqtOC6iikIhihc4mc2Anp1WdAJASu
vshBmBAXqKq+/hOw+WLFzKEAXMfCnpBhPKVgBasOXJWrOewveqxBLouqahTYQsPHv5mv0tDwkcjD
gg0GmkO12Bv5xy80jNBFw/WqKH/qPmN80a4cl+4HcQmOv3KOloe4Js1oICemuOVSYNPy6SreNeNW
KH2LUFntuDunxqI3yu/Vs7DXLwsJwwxqDde6N4DIAPGzH+PzCYjHWteL8I+Brbw2TYUg9ufQqk8v
xlwdQ+xiTS2MjpyV2CSfBykS3QsAvmlb/tGhfJUqQGLUGcI0JrR6AneF3Ae8d9nfzRTMO/cS4Pbf
WdHHjNyGFPOM0Na9Dd4xhXSGTbDTRKuLgP+2B+GWZH5Ipk2e+lXwEMZY0Z6gFE2bdeyStY8D4AEg
x9UcwOaXpyp8iHEOoaZjdKrdvVhMx2YrJGl6XWTilSXesmQjSFbFCbL5obkAmZvx+ysp5JMM/QTS
94ifVRvkDZCBd1qm5XhzyAl/Cg+d7TwuwfFcM5Ix51VIQdeI67PtHdt7+1bGFzI/9YZdnMJ3tNtb
L5vGs8YGsKBmRfo7sp88VHIQDWLJXJBa5GfntEeJlPgsg0nz8tFCDhYiiNDdU1/Xwd5rmudEPQVT
w5NfVIyuDYk10vroI3mgr0AkkuszB12PAVEig/EmB6MH8eIS0Ouv5ac8kxtK1b1PAHoqTuuiOyX2
Rqzv0dBKDPDVEAUb4cL+T2KH19RskgOtmpBvxJUxYQnkCJypsnSRliVPVw9Tb2eGWToDtcGTr7vU
8KM9DaXATvDqs1TT6TlChB68QkB2lMYvO8sPyGAPVOwn8uL6ppscpH3hptZBPpRU4XrXaSeRCkuA
YbmKzqe2BG+KTssK8doCF/xAap4kqkLslD58PhQAvp+XOnDYOxcUiz/c2ImyQkSdAPhaOK+il46P
D/BOyJPqkK1KrTsgnFXwibAOX5LfvBpjAqvotVkKvOkhq4n58JZ5GYqxWXPX4T48WYhift6UEB72
+m3z3Ww+Qf64+xjFbMq3CFdem7tu8l32iGDAKOTO6o33sNr1JY9C9eaJYykbywkQHBtuIC0wyUhl
X4yinf+0wCCLDwo8Vv386IRROimS3llnUmC9ZAFn7TfpPzcJy6LyoM8vYk9x4lJ6nCrF/cucXQ96
vTRMNzbSC1H+T4NaYhfC4jEX5MGVhhflKgIa4WFtf1qkPidZjUyRqNFdPBEjhbkur4wnE2cbDl5D
VRWUiM0sLQCYmPYlg5Oo0HF9XvGHkIOpo4HZ4DG129ynBhqoXEHq3y+7EnPX0jTBatz7rfFyYkCs
8olGyibHAzH4v3bMPIc72WE+9T2uA/JMPmvZRWptyPkurfizI92BOiwo+8bHGI5d4anYOx9KTPz/
CsATL/sxQbLt0N2wzf9zwWZ91x9OnaBdxWHWInjkAMImYUEmNl4Rdyz1IE0dTlPZlkO2SaA24fGr
aPXipKTUWJ8+dtgBfh3xeJwdanP3wr4XgaSaqdI8TSYtRYcXPJlX0QpGcxqtBefT3/uyApOq/pb1
BWM/ePk1y0n6f99ZEMaL5Nbkzy73PHstwHRQP7upkzcoYqg3nn4Bl2XJq4gBmsV8P76oKAxxYkbO
oigNEpxQYZvP4rDI88+RsEJW3+dPsp8ne4qAdCGRGYl8+PFHBLj1SuHgKsMtas340te/VQP3ZosJ
RKy5aOdYf+h+uHFqSUb0LSRaK8KIZn08ZOyFcOV8hsbSwFfrPYTD+xRuMTmvvdfhhdgINBlL8wxt
TFuNg4Jwb/QN8p7ZbEqLr5F4NLw0BowIYv7AfoF81O3r91buP4aJPIMptgWHcoVTIYTlLCzp2ItA
wNirkvvYgqWmeT3UcdwXwcE8ltAbv5JqgZi6q5oi9BWCBJTnxLY4f4DXmEDbYN7bT7xC7C8FJT/X
9nhTJHoMiQb1rB3MtvJblwJE6snoUVuDEZhr/g5SseYBZUtcOWJSPFn+ym7Q4WAjP+EdJXP20JUG
glEHycp83neXG+E+eLBmmrLe7Z3NFGBEg2AzltfiMz+GBVMoAnr69IoKn4LFCcAfLCD3iticovtO
0DxkYDndp2jFkzz3V0+Ig3jWSlsNpHWu0wxKWFjP+F2DNzzUDN0ZdRRcIAWAbTQSPaqke+kahWu9
GqZLvCMEhb5BihBY4vKmchY7IaH+G4DcxNV3XTR1jCDVGQ/JEKHn1RWfPnkk4KmVso1VjcymMo0n
6YrGSZfHLkrEIrCbccuic2TamW2UZjPxRPgT8ri5zBKcjYu9/qS/cxITfX3iFd6MuYnGprjIxXMf
2TefHysTNnh+Ke8Se1bP/X3uSxOSStr7192wqWzqP/qCJTLoMgBprzfgYhccYqs9IO7mW0bTDcpD
z23JFc7u7fPAPvJYqMbiblWpke2GUPRHWn7GRR1pX12c+ItDjVizST08t79rRlFZPb5xnO1XeMZT
mtyWQQCygFWFQgSNY8qAyXq4NjuhIiTgT73VquWwQF8IkhcpT7S/2iM02Jkh5jn3aLYYq+oi0gpz
Nn/nADW1J1Gz68FFemQV0/44oRoWV/XdE9n8bzjlF9Rr2Qe0hYm42dheWIyN/D+hN0vCZroyy2WV
RC+Zzk/8oXB133al2rSCqiOpnVbxI09WZdao5tlpRof9hrGwHyLx8JyixdJobEDGGv0Gy2OOpihB
LzJd3KR/cfEgGnkAkR1g3x5xdWwGaCD4WlPHySM1wShT8WbrSqemBOx57bzqgbwcGYTrnywymgAN
S2oOtwrCLNldbw8K0C0fbeM9NEwReU9/CHfrhoASuKDIW+MNMXnCY7tAva7EXgBzBBJZkb8lAhig
8mt9HjtcTj5Z/QwvQbsnWslM4xFGlxI6V+wGaYKO7yYhNJT7vKV0riiEn/qhk/jXvGq/uKtwb8Q9
Kk/5g95RPmUggAM32iKBPRn84GsaQIVyxhNbmu6ULLzOF7Ub7xeL+Bttw035hkJwvM4UaaN8G/cK
QtQDH1XEzkAjypBwpRuEmIs0dzT78WBO5nABYVTrwMk8IKv4AIXi9dLhxfHDcwhBBCeu8dpYpZ4q
zZU40VzSlMc0YBp2miKDDmojEeLlZfb1Hprbwy7Bxz6sohhD5qd/+vtuC2jEwSmn9gs/+FaBw6vB
Au2E0Wr3CU7lE3TXp4l+TH1Dnc4yE3IlsZhYSkQ1Nq1+SJalPwIW2Wsq6yjJ7ZPEIG/V09WPFqqI
h1ZVXjzvF383lbXo6lEGFb8yf6HncruKTm8QrhH0YHyB2o+tsdlTicH4zzNCIMwwb+TkH4tMvM1R
jh/TnVhwTl/rqFUsTC/jfoW2BhMCAoVzIcIFTz6Dj4iJBBhBC5OlZ8uV+m6eJVjR94ofN1q7ZRMw
aWJyduNFBBjRlITeAAhXKi9l5Td7kwFJ4Fr6vDcsrvHI48wJiLdil0/+miicP5PLvwKJ9vHyXKM5
jDxActWpZBpbjf2IcgKBKu2BhXCLbR4apdeaRTmyC0ds+khMBdJqfGjmsRPx4XCyXQyEk5YVSCcH
zdI6pjRunOY5YQ4lx2MGIcLofFjsqE7mU+mtLnN1TuiG0jWfetAkA+wHTqvW1o3FJurxUMZHqMrM
01fRcGxJTrqPS2GmDiMYHknKccYkh3qog44/tfsIZJb+bSjCHCveFtlOdQmNwoNC2aGMt4zN699X
mDITl+3RN78QUVJBi/3EXSBfvWEWPLvMuq8OEhgJk7Kgk1cMit8DeGhXyBXh1OD5BWnw+1MCU1u+
nkyHvQwEehXYs7MW/GeKp32IpUYMMJrdNRAtEswCvC/3pk/ZejDju89XNfaTp9rio9rYl/6EO6Qc
P9preuU2fvbJ6lPCgRdhOGUvERkaJwcfqGpNOAgOxFvRZYSZLaUsjt6SJ1DBIeYRmKoHTDtS2vak
jJqbVujJjC5rlB0Q9qlqsLbSjki1plm4Jjen0ZsDJ/bSB0cWywnr6jNqp2/qUDdehnoaM3wrVKJr
nkSB2bpIKvDnAr/NK9jTQXgBqMvcjVz0jMEDEdZjUuPMtT770uJFls+GyUoCyRYbf9NNZM0V3kTf
G3gNwHQlZkT1ytVC7iYigN0XeBmO30jQ5ZqUvrB2MjYVZdmS+ayWxzpkVgrjJMyfoe7Xp39zX1aL
b21Di8nSmCm+KEr+tWp87ICko/LXWs0Q+IdXUmwgirfPHZ97yhHgSLps6c4RUaiGx4s9F3tvyZeA
7KnxNV/KKZU78jNouhM1jlKwNrYnQNG8/ClTCZUqzSJHoSG4+bBnRQs9yvPwmhmmMdR400L1Ptch
LatbSr8mZIDql4iSHBz7ibzGNd4F6twlOOQTs9mGPGCJDcdnRAze2YApB+qSdJltddf1ZsBxYdt9
S0Fpid1h2cmEB3/v53qLpaSA/jB8+SccVk/CiSmJVvysW+vCoQMD0THDseEz+GwC/gEeVuGdmUd6
7Ll3Q3XDl/ZzFqJK2SqrM1tbHHhboLE0D2X6VneOgjBqawdf1c+FmG9JZS3EZc7G/Q6QfroDhdIE
LX+hNOua7NeZ11o+rZCamRa4hOqcZtt9hFllkkWx+zH4EXvxZ6o1h7duCKKN78U5RTu/Oi1RHIFL
zkPCQ4R962Hwp3U5nCtQf6yFTTivemBEE0zxD0RHH0OIRywLjOy/g/gjEgrz+N3CVMqz02yCos8N
bS4budyXYiKBEeFuXcKuyN1WpfLwYa5cSo+/jyByKSchmT0jowO/nj/r6GmQ/2ux1Qj+LBbuEfAw
rCmtfYtoKFeBGG//HScOoPJ96n5M17+q4UW/bVJTxNKCtf23MhhZS4Qqm1Sq0nS8hRLOFAhqZs7W
8BX5piiUsFjmNqZq0LKxnZ0yuHGoZygkceSFofPdlkFBaqD2hNypWVLHWw+kUT1sqtFp8+cacteL
7jsB2XcIYuVMo7Qv/uDUKO1Q9DqZ90bSthmIFMj8xe40I0clAWBdjysHyW7bMwHpxtLD2que1LVw
98SUy39LV+AKlyEtJxQ+qF02JN06v7w3jE8Jgs08vq5PANg/CDAplvJrMz5+O2d/mQi+ZaF/SOQx
U7FPQISRlXu8wDm1jtn8bNb3c8mgQRcsaP48QrrJRzrVIq4N6iOHTKzOZBuGH7OBu5Ge/OMXiYAH
ePyo7cy5FLBmZra3kmN8fbLol/jkIwQletc+/w5ZcY2TfLldIApE2lqMs/mCFYAe2Wj8CRACeadU
S/kHUFQ8gw48qlHy5yajOkstu+K+/9KMFPPuY1yHW54plCKJDmehT2dVNZiC/FaaCd1FhVtbJ7XX
dDE95MrzGm9AWBXkBJ6NvM+tszsmBvKzEU8yihFYXTv6qhAHLRiK/NzoqvSt/oxjb2UunU36LtzO
cqHx0gyn7+PAoBcrOkL2vkupFvWRhaqTNxHWXvNhRBOrPDfiuGQim4HxPsOWRRKb8t0d5h+ybuM8
ii/AA3PyPIlatRqdEG2+WjxyA1/5P7y5w1NHqFkiuc13wdZts7JgKCv9m14zgZbJP5v+gCG3XdVl
30geTBJts4uC9nXs7cVbq5VsDv68EfS6Ei33G64bw1BY8M6EHiVVHjJenZ4N6dGXul1U9qjzry7D
wieaeyK28KWaYbYJs/uc7n4ohs1jQEbM2noXpPwEXly4sxJaPxqg7KFbsPsZaeDY9zABtc7phuN2
o4eeI2E6dgPtdBjeQzy6uxzluN6FH0xTL5No4iZZYQyUFgzKsPJ7rPiwbWC8S+928QYrZEB4F15P
8sGU0/arncswqwgycMv94Zvrj4dPULTZfBPzkkwDGOLVtbHN6Muhi895wnA2VsG0C8SnD7ESsMXP
+rEgtlxnM6wH1IKLuE67Hn+8xkrFEC/HOn0WUhVObmrc816guSK5Mb8UXweuCuUY6PfpSAb3+Wfy
8hY6nDBE678Kike6425EM3d1dUP9mlZlSfh2D9J2NZ06XvxHgnD8g/VP83LlXXIp93ji1dycoyyx
4QZxFm5v4NXUclOBXseyX2QMmcPUaEn1TTl3Nh+QdyOBkOdBQMu+Cso+KE7aR7ywIYfaJxI+RlL/
4J5+/Ko3NNyipWmRbwkdoW9k0oSty2Lpsc+62T6pko5Ad970e/Fa1IBdM1DPHwzHxdOUEz0dfOfu
0lWUYRX89c7Iz0ID0W2W0ZRM964InuqwiVjua63771ImF/YjKb1KeuRo+1uA1A9fIKvAH8w9uMUH
p+jUNR8pmSxa0OqBgIAxOGtMKMTm0hOPiAVewmwIvUACFLFbV6pnEAVHMaBQLpNed/YZXzC3/8Wi
baFxamSJtOnBGy3d/5y1X0oEvQMmB5ldNxZ6ng7e/Omy1w0JnJNqtzr16Sc5ICtHZuK+t7Zq0ohl
Jf7GLQf2ORmSWXoPuoaBWeYI5igu5K/QYEhDEipLL88Sai1yyuSg/XL7tKSBl6UOZ3JrtQFlhycM
7WMErc5R3KOqj+HK48002rRnkMPKESyKoIPfHh2hpWcoJjwu4qqh7QIJC30o1EGybJNfim59WLrU
NTXILxUIWHc8M1ut2M7qlhJg3zdxE2WSXP7jJu3QRG+dgziLVUpWCgeEMnCIQUWh9xS66LJDIKdA
4ECFUdEVxJGG4hmd/5nWcKY7DFv7A/oqgXGKvWIHqJDmWbuDtmIIuoY2ccoIhAJh1OeNexf8ayNg
TjhH8WNeFI+6llvkRF1AMER41ZLqxAi+7fXZPAD6Cqrq4OTg4/MV1X3vJVk8grnToDy5vAXt0Zw0
lIh300cSMOjWxGcjQr+1blK3oBcWtHizvSQ67Q2cVfcQ1O4UOwxB0lNZhDG6CyzsplaEeH+YFZAK
AmEqYlsPihuUixRCmeLf9PnR+A7QYH9vPgcHWwViWErhVMFJ5z1oIAJBZyI2uBal1jQya4nlVzEr
Rm+0nbsw+AhRVJfpdwhhiR8uEMb0CuJRwoZc8zduW+5O2a7PQ3Yc6j3BvzsrYgWRtfSucdOMdp+X
7Z+gkuVfvpS+Hcp4s5AuqwKJvetpOQrVrylsenK0B5LzYSLCll9zPb95TqCESnRNY6kwwE3Dnsr9
F8pYa6X1P0EcxntPJv1HV1l+/paem0d15ctZE7AeD6T4bjQR0BXbojElTaRKYfhXNJl/TCtFMyxW
cuZA0F49dlXa8P2vIefIWOMrtwv2sT0nuZnzWrRsIEA893NshFYaIy67P58y2rIt7A9Sh0AqyR2F
9waJTgRtIDX/RB+F1L2QVUYtIcuUZWLuxEWtu5jjDqZnlHVMG1CUsOKTdKpBtcGXcKoSZwmuJx1A
AqOROip7iXc/GIiDp6t0R4+k8NktKI/ql5B8e84imVZMCPrEI1ZeCxsJdBBO+Pk3wt8/Sa1b+rb3
hUSydjlwOhDnO+ZPaZ4+sL6tp/jRTz5VOxhdCioRsOmn712awezyJM/tbEPeMLFxRUoArvTaT8z3
uQSGXzDKabHMXBll4JkPllXyQQhvsmhO8FawsHDuMdu1Z86zPf60pfmqVSOK5BDM45WQSbhdQUYg
bTDS39h+aM7uxD9MYbTxNpYrDdX95/+jpeE3uXYXtsjJUxckW2tet0DIT1QnUzUiWB4j6MCP7g4r
KgL8zTat0d6H836fhE8ODzWhOa6b+XbyWERtWrq8UX773uEbNd56cmq3exDIhYw/ekZYOugpfdaL
uEiZchd8f0Uy5AfLAoac//F0Ae+nuD1joDYuml6tPhOFlAaUzCL+mOP0ZkWIWbGiUrSZP54eClpV
l5txol7X9yIwQefySO076woMv6LtWv8qaLsb2GyeJ9Whmp3JdbZIgyih8RCpXaY96IsY1zlidQhd
sibjqaI7XzoXqmCXPjIcRW4faBTyGPASX0RqCT3tWLv9ijhIKqMir2G/ojEdmXW6UFWVevy+gd74
pB/V33f3DvxPJnHCohlhSiX85Til25k6EgOPf2tkM/HDguYP8s/I6+A6SrBCf3fcHGTlD4krBCto
/nw5hj/PRCoWvydQ+k1BLTZkKhrZ3vcuEr3O1gMSmv0435YjJ/H8nzfqiCHTla14XQAZJnx83O9K
fpnXzcFpCkzoR85Qvih5FUiGGvl2bO2uBO/jwATtANjt/2RR+6KzKwx/t4ZuAyfB3/jptGeA3t6f
ReN3SCqZUuAY3TD6jzy79X6U0ZAHetcNKkQfevmaEaSKPQYXyuw69pojXUKvr7xviRTYrSof7PSb
Bp7k+gL7Q9ymvC0Txm5qMTysw+/aSB8vVLByr4p38+Ric7YzeaDBGuthEnYLm3tz9Jiw7DLNBoXY
2BC2y6SIlsK6JLLICk592KYaZocQtzqROLC5bNEizRkK1/GG+Yb6msbb2ojFxA0dUVSzb5itMMDi
aeHkqs61vQYriy5mq+HZ3JeShu1ILg9EW/pVo4y92+V4zN1Kegsq9lVKPRiDrRrDVhk+tRgkas66
cQgxTwqCQ70xBkcxAf4hb1456A5+yESjfZmOUNhPUAmZgdTzNWjVmzCIGHhYZFQBWr5xoy/+EHNz
0ECJB92ktInMsADNKMCHG6oTUQmitDmPPLJSxC+vfFBQxjzI9AYu92gTn9Vb9IKPnbtbdkYrju4C
7+4ij8nl48Ik1JjgLwH+DyP33or1VJ0n5JyCeV9nsEFbbKQRORm2aFkQIhwUooxkGcIfvKWT7WXD
JX6Wbn1MhLdRETuPzYYJ90OBlTiJc3RuhGGiiwfjj8nd8DUFlnw/rb+Fa2vEZzkiaMIFG5mG33tZ
RIpAiid2q0y7N2LUT53KjOr/wsBQfIlr0+71xjlMgE23GCcxrFrrSdUn/1EojX4dV7RnZKR4aHIo
kktprTxmDyTC7SLjZDenplqjP7aAUR0dVpaEn3Ik1SepLFgnhbU536gjvlznLlHQJdmrB3E3WQx3
gn12HrZvsJR0l9ppImtxWGVHGokuzlhvH8o83MxQSivG0i6dpZzQWK1hkGjLLhXpBKBKDYNejL2z
XyXxO8MPuPP2UE9rqX/wFJfRoPFBp7T4bCF7YyoU0Oi00/UzpjpwdXbS7EzC302kHPGnIvliYulO
KD7Vxhb/SMYOUFpiJj1/l36gOxibBRgV8eCBQO+vTYCDSJz26AsU6axbR3/+ypBPiu6QRvZkFKai
rJCYVoIkV0JyuUsLVAvwPVq0v2JSA05TkgZiX0mqwX8VIv/GyiBPNSDaX2QrKt6DASVOJdnaNXl3
MCDoKtU8HoZOkNQK7XklNjpS+ELYx9AE1w50xsHemmXElfW+MFo8rjRzrbrnLBNp/kYqKTacUhKy
J572ICeUxxx4//nKOaA/bw/qEov7XxOlK4vQG51q2CyuJIPcGEmME7X58PKTNjZstcnOMcJ5gGXq
1HsFyu04XIUTWHKIam+zcgxYbVvXP5OAcjuMb0R6JAxQyysyB+wE/5vDmODou0m5XAilrWlLFAxg
eMSgdUlWI9YX2XLKa0fUC0Xw53hDrMYzsYjxMBkRtOIoOASn31VxAKFV2DsZnE0U1VPZs2vO3kay
kDOw/zHVjoug/j+6zw2B1X0McWYJ5Wx/0tX/kV0+cIrKztQ0zTyO4zP/8zgXJZbwD6xS2dOIBYrA
9TZS2kbwA/ze29lO8EzTjObf21frbJDANfvPlbW85QWoYHwpHiF78FjZKx7qHS70uXOiUFWe4L5g
pZr7S2ckxbZGKxi0NtiJzGv+co/5JVag23MrjuPMRMSw42Xs9PsCwKvqSaD0wFd88q1NLYTpJiA8
tEpstrHUYOCRRLYx3F+unBX6BbaNUP0/mnaNe5EPJ54mH8dA8Evl+hQxW0UDa3GvYaaUEE9+1fqq
QxaeHc9qOqzAf/dPHcYhwmyrFcjk7CKfVSklFPegDhvocwp/hplla37dZIEVwCmsOtaGCcS2WqRX
4ff8mpJaZILDnHY6LeoufmhnAynkC9Dsf8Mh4HRAvgE+Mwcvq9+z7TkK8+KPBzYpAg/XF2uGTP4t
W6wGR0nwdeizudXn4KTwHACk3XYDDAKJkwzPhg4JfotDb+ocnzL8yuJka7+8P5HwoDHqY+NRalh6
UHEkbdAAgcqE/UsaH6kL7gh0AONqI7Xb/yUTyLsTT5/EoljMQZgzOankuFnTMQP2uybbksBaeuTz
V+QqXFZePH+lYcVcvMB/6jWP2marpUou9APO4lzIPRc6S5xfapq9eJxYkdAS1of07/J8B1qqau8O
/m1PX488J+JQOK5jvTpUn3NdVe9ipupu4uxqF2l+4TFs349o+F3+udEVX2KcAlKxT17AYM90ZukE
6O8i+52TW3H/LpdfU7Zwdi/YxT9OU+J/nDgN3BJfIHnGGS3GERjuTaptFsgfJl/1oTceU1YvdBnk
pzAA1n6xtwQSiYh6NvLl1WQ6fCpR/T1erIS1J1EYjTISNyA3ETk04PsYq0unnCRqqgU/2WD2WdLO
8/Pp3NqAvAlBhU7HTeZHdYgsPac9BRGVMyXdi/i5xKh/BmLwckhpst+vbn2qiNe/p1AlQFCGmTnL
5BjToLG88khEsPZ79H85zMI1JelAyshTt7zkTcBO3PIRmqvIUE3UXWi75MrLAuE8nmAFEhg/HlKS
QSOk7GPUJ5Wo5YHLI0vPJA0iAejETjTHCGg8M/CYH9xHmDZu2snPZz13HWnFfS0WzzG8UQOxFxkc
9pT91K/Xk47MqmjBnSXCZ3ijKWem+phapi87Q+JPMP3dY8K/1ik+ilKAz/MQ2cYwSNifB+TdTt7u
ZkZfTqsN4y/uG6DntYShbwlItxk9f3m7aA1bp+8WCzZ1FOod6bp61Im19iFprSBMaeg0b1F4dOyE
YCxmif12s9zqEJ0xaA/yCZKv3PzhSbVcB3ijZ1Zm0K0ImEcY4y4TqC4TLI4BVmj3fDPvJQ09fy3Y
BRxxZBWPI3UDxYR4vs8pcogSvuobg5oSK6z553NycOsfj5hC9euTgdRMb1q/ynqrFQFd1ewCZGna
XvcpxA0B85iv5xphr4UA8J+Mccc2VDgwar6A2ijXmWoLXg9GQv73s0VQ8zBANZq6U+T2YLflBquq
dM9LZb67f4SMZMm+X+aCkJ5rL4xChEjkrpPkPyAqgluAFaIE7JdnXn/+3JOCu+dLUL7zezCxUVvl
ar0IEH+eSeVPKWtHQtO//tDHZOxR7k6uELrq+q37xggvc/2nUFZBZYR3kj+tjSGP53vNMcYHDjl7
sbWkD5Ix2HWRkyA5iD3/As34o7ci92NTgXd12EhO/s2jTq9wO7WUGosWYzBoObb0oN50E+Az2Q0h
8Xx/2iTaCbh5kDQN1uzt9XqJc3SqFUZBg0+I55+U1M5C1XDdsr6Lv8npML+8AkBVHzgAuobYfNb2
p5f6aTscZbvek1YfFVhtyXojUc4zLwKsL0kopNPvYOhhSQU4M6ZVrOePfdhDCrVaWVYEF3yavs7b
9GJnciGzEiZPwSMlw5TYiDi+AT6zmnK6AHZy4BEHRP+BkmIWJO6ifPhvCh1KNTQ8QDkDXRAypHZM
rko1/izo5G7WhDlIXX7Ilk0t+q6rRhvqVba+xvfjXW6qZFpRkvt5wKHrjine0w/ateujT41tVxKp
AwfDyb/+i7E0yK8vkGHMHws9RBdmBUNJZDhnkD6yV4h/3+EFCkX8cMuXw2vbnnN8Qiahn9bpcoVE
7PyH/electJeg4aZoGrkxralkEde6Dsc92QHj9G/u3xr45LjyFEVquDQ/rhpj2a91xF0iRjE1txd
DhQvURgMBxDpu1XhBWmh7SQ42WqK6LM+vJ53VmwdWEOywfgY960XsnMhj8wUeuGCmZpEtidm1u16
v+IRnOrVLGCqYREWiK7Dkpax72vkRdV95Pih1yQ+6yqf7mk5gizfMsfhy2CJo0+4Kp3wehBh0De3
H65GtOtAeuxw6gfLVNic6RCnmdH3RMJEhNcys9fhAjY5E6XpkhwP60684DC9DRHzlo6tA8TSisAR
BjgChfCctM6NJLHEwGVp96hp6WiYURdSBqDdsm1Fd1LVNZ4Ga5rZtVpFjLHsvV7188P8x/owCoNF
JDkTsVh1Ab5w11QNJWrVieT8NswdSHn+w8Wgt4ca4IznPY9c6rkmnU7fulj8YD/6U/mFMoiLjn2R
nABekGssocCBT3T8lgl9EY2G4NQgHobJ+DTuGuCrQFd+/yngmsK1wKgmESY5XLIQbTdhFom05YBU
fw1erh+hcAARQ/zY+y9ype3bF70Y+DcvNW2GoS/hqXaG83F0meaN2hTDu/WYA1jrRHN76dzi0IQ+
tMdAe+vKbv4waVlcF2pYKfhzn1T1hKKlpP4EUahQdPe+pKM67Uf0W7aa48zI3PphY0MDZjgTfwhW
fgW/1B2gwKyuxrXRmji6gETbT/WpT1Bw0QOG63A3ks+L3dOa5Ujsb+zWVDnHT0QAWx5QoJlqvpYr
a2Vu4uCw6hIs8nsvroOWvD2LEhqCDj4OqjG5h2+rLi44+zLZ9m6s3vzNLEYFOj8wW7Qb4seka+Wg
4iMMMKj8jBGrQFsW+e2rlRc1NLdFmICJ2ACEjHiPH5JwiBl1QB39yWRyihVNpeKLJ2YC2QZmTDkS
jYBDEZGTdexlXA8X4XDlqFcNGZr+ocQV0+yV+wWLDlIeX4HhP7GU6crgeRFs19tUr7e77KhFkoSf
Uvo+zWcSAllCEbkQZD7pPg72wD+4ha6BRDgo48zV6Vf2e/pmubm5fc/53hMpmLRGp3H+cdmaf40i
xKFNPE/+AhDCmFrHl+zDJ4wGgMReOj3GVcPTYTPQ7r1dLId0AHIhD6l4STbwQM6BEGQ21Fm4b88t
GIxlI9jsXJDPa7xYlnZGWPoP2Iay8i1Xs7UcxndLqXGefVlkJLmWMzyAMDwk7yD/Pu3KkcwjZk4j
uzi57eZzrfRSnJPmO50XL0Og4dAyi/C8kMJjuqs9O/KxdTyIlwVtI44Vo0tbMQtke7JANNr/TiDl
5fCY/Y4+SH9CnlP8LKyxJY/GpklCQf6ArHag7PBlcrRRQbhhGyeq1/F0pmhTcAizAbgciOdbL29i
q3eoVrhcXsY4sq0qwaFIDJ45B2oxq5nlj3wJ84jDfxAVztgcUKACP4z+AH6/vZXUf27+DGwWIMwU
Gku+ZmnHFWMXgRRArZmsoPkc4YLDM5RyGnro+8VAULV5VuD3Lv1Wp0Z2V0WhEZzeCevgnxASwLcY
hAKhZvGtySS6ZZWJEHOKBhuOgdygjV7rQU0nStzM1EhVK8o6sgQz+i7lwb8g4/jH8Ii3zmDyo2PX
PJf49me8Hi5DXqjcetZoh6JMQUb3/P1elhJ46uMVe/rgX5ajr2CDy7emn6j7E+hDVyxYFqFv3LvV
sQdQHjT8hmbp1WVyBL36c5lcn/Y3llMdYCRVdKknTwiYgC1+Y4AhzM3eYlvdmd7D7IdORB9v12Xv
FuLRieLOTsi7v4glh4a6g201ak2N3brDf8zcy/9b3sd4Y/voyDsaiM1mo70ELRy79h1BZBa+w/ee
xOx0tiVcdgvOa25SPbrnZanvJTsItRW96XArJiB2m1QXG/ezL8KxMdk5S0Qviknb9mq45G9Do4P4
xjdnOAoFVGf7NbrI1pMULDR/uFddJtJimli/x6wTHWEJ6QfvSdIwmAmTYo2MJqEiVdhkW8Qzt+b0
BBNkNmFxnP0xLsmCVhNJXIzqJ+BnrPt+IEJbMyJG7gwa0dhbSXOtkRoD/FEXbonSNxOg/Kkbv2YK
Iv3UL6Z86aNKyfz9T81cyTd440wN2IfV/emll2MFsAycccOU1Y7WyR73tfuUhNzpsT3mYE6gPn7x
MsyUJRDt8IS5ettWf22bJznlWYkU6/25Q9vXLNY7QDpf2y3shcki0uCG+LrDrRmhhfsC8MJElX4r
xe+TKmAs+gHSY4PSL7LHoB6GY6qBGvnELXaRambKcZIiByC6PeZM4yoq2D8hlJ8LlKNhK5kFMKJ0
+rZ54vaLQPdIivt3i8IR0eYipcr6Ma5FetLZMLOT+9wWz/A/SxOtfRRz/V2EQZa76wTi1Im1Dg2c
8b0je2tc+XQaxeNFGziElqXXNQWJ2uAlQtSm4bqoJP9chJ2DzxaJd0PlgVhrM1sCNe04xicdzahs
8403cCc4QteZ7dhW4UDZU5tLY6UlEPN12yTQGMGu5IH6LodeyadGCX3ImMh4oYkZG4gT8Y7ygSfB
SnKMB+h21R2MmVfZObqROKJnzu9DSK2ZhIDzgq5pThw3E9cUQpjA2m/Qfd4s/Taii5toZVBQWcMe
+b8gsI76rFdasj5jMeVm7YRqibjw+sKtZALaDMNv/w/JjiEiZgeLrdpRPE/2+8iykGzUCjpe45N/
da2S9Yz8yjRWetIQpj2MYvZFoNwssZbJTZEX2Lw99ALdNwnjxP6AkKvLhhOnpru+8S6WmhTvjWUA
3z5/jWNbehDZXcqHfQiKFI1L3EoQ4Vu7c8VInotkZMr5OKHETuR9jRRq+V2R+qroKNGX+sVr6KPT
EvPhlTiFm05dOjFxsD7UcSJcWeRyGzCBBwsZGGlLNszh0U1Su7lr9mytcpGP1rb23ZjfmRkyldM8
IJbIbcqaWSG+te5XELhcJRg5K/KgGr2ogXadU75Xs9RSQ/vCEKMkB8JshR2i+O8Tf0+pvfkJjNLP
eZllqtEBP66GqM99VFNLTpoxmIpqOGU/0c8QZCvAm+ts4ZHfvz6/zCSV20hBuzoB62r2ZbsN4pn9
ynsVqoQ/ESax+89iaffkVqoYF8D3t0FjDBRC28t79yeDzLRkSl1U7pJsq3vmZj4pMu+TTyIJUYtA
xHprtwX5N0CJNkhT6gkPpI5z4PlWgnc6NoIqnEpoLl2U7sctOrbofrZL2gEbSXHxP2V4QnQVbAu2
KttVSVOcdPLTKU+rtJhaP3eK24XFSiHeKLjw1NMeCkYnzb/McBK3tSbzDZpfxeLbcGK2nefaKGYj
iwLtNQ10TzXzsPiR8kyyhpXWips5cC0zN8KRGGoVA1UREGSQihPeHRNCU8st4KzNLlQzTcKhFPWR
T9yKXHqAimF37KpBP5Wd/eip/fWdSqmNqA40ZndfW+zi5ffjDERkIHHvD7QB27/jQ4Ug3ykjpogi
Iv/yMTpDP4tg5XmxK8oNooIHXTb/2YlBfw82+Vg3Fi/ForiJK3+QzD1vvHWYQPK9Z5lHOG7vcEBp
rGad/0VXDR0ib0uVZVPuZQGzlOrjlsY5SICQNBA3BnOrfQYkRFHT4vMMpykwIAuGVs81yWhhAsF3
hDoLInYSppJBDsxbiOSY50R4X4Ea5gGWkZ+0V07vpm0asWgNaZDDfAvg0TwsbjSJxAc+aYvDphs2
4M8ksEE241IcpSGmhfcPlvRXgm3HSJDuAvR1NK9dCP6Me2a3/MY/tyUy4Tme27IQ5tQ2bmk0B5nE
x/kCG2jh0DiQf9xjL64u7B9N0MK2dxdHll6AXosfEPhz7eM3IsoTQmapq11kg+5N5SldiLchcFY/
I0mOiE1RdroCz7G7kNN8Q5soXUMx9Kp1I5CMt9P8tKrOL1SzbbXYUwvOUK+UrEe69jRBvt3s69Id
aQOBEZKXO+zanQWcpt/DNfc3U3x5DwhKTIbGTKjCbqaDBbqTUJq+sQcJ1XW0s+yAh/+8q8Jyp+AG
y3dnTwgQ6/Hb4WakpGv/3G9QJPx3F4Pn9ndstHjwrKquR+QK+9jITI0PZ5f/wkOJrWDoVBYnvk0Y
hBilXXHMIijMM74gGnFDFRMzXgo49TS7YEPZc5QfXIBPgCGuHNnJ5mSMH7RKqroqyZDSU7Ty56zi
LCRjJm1d5eu8b+QctOG8m9msCe651+1snyeBxtQfDhWGrgNK5BqA27QN5G05/JrrByM0WZJGAJjz
G7Z/t1XR9B9fglqASAOaLsh5Gq/jJHV5Q4vMmY51Y0w19El114snIQy9neGqGLpGZYm9a04f40Hk
++xC8C6/CGToRsYpfAUUsWegETF3jC94MAjHz13WXgBr+MgRbcLqpH4h+ldtfdBzNTmsmCXa6h30
wUUxTWjtqyw9Nv43KnOoO6g/+shxjKqVQaDljBp4dBl3qUA8aVyEDn4p5ASDqqqRLr1KSPqlETUx
WUNRoVdpUe9+LwyuNfdRiQhqpJq/XqjgeLwSddMd0sXHSG5+CBF8pu8eudx9gtcVlir3wRKLI10p
nXiODbwBzz5nxWaLi8YU3o0uXYhCSnkWQu9xq4rMS2wnKDDdpPZzXl6NzevthAf9N3PtHKH7w+cP
hC5UdY+1+NbGWuV3N+e6TKoKvjzQgAl0qXAptXKuTJcp1xAgWaeTb+b5FR6bR+hrRhLjwkKuTSRk
SNER13Qaw19+fYfu5EXR4KDIs+OenBaG4okpZqFHcWPhRM1O+byB9YuEHQcC3PoRXSU+36MeYNhX
mYmVbqHaL4Rt8ihQiRBA3K366UxlITvxfLTqYLBxsF+UG0/09FDllhTz/x9ChftbrSuY4GYDnWAO
BKE6A3UhDVommvguEXg388+TgRtZQ/u0wG5DxA6NY1Oej0MKUXNGHdVAw4KvjK2N1pPJ8CXmNBdy
0O//QJf9/UpYH8NXxxu2aRzZM7PgiBcViu5X84Q0376nbfNVBVbCcNTAr8LrkpG4ZTYbxxBdgEE/
0RN3HVjybzevEuEXBOO+bk4GeOCLu0zxW1xLUcId4IBOEHcheVldihK4y2sXhCvfK54W+inO1Ww2
OhbXhoY5bI6MWPP8QCtKCaAWB1K0fucobNyGUFJsYtYn1+qpWBxTKPGmKmU85KiqZfkJokCFC696
0iAkkiweF1uc1VdWo1Cdu/oTNjuTCu0CpmV2tZSLIWgMR+LJafOcYQ8B8tPF/H3CB1OP4AVCfbP/
t4Ii1QA1ELBJbXD5KWVNx003i29KQwl9TtIYS/N5z9sf6p/Exys3FYUnBV0MM6mPupYrgTVzJ2fI
15ynmeasy9Hd7gJPS1waWZxdBZw6cwTWYm+J78J2bgc0v+usUDoLZ2lsHX/XTEVplBUX8vRiNOKz
s7lMsLgGCav7RL5SEAL3mlBqgo/997g9JGhMrIlqQzD+JbsKIEIlUE+BTqUXkss3AQVgorJyqjzu
yK3HXjlloXy0Qi1M6/bKOkHPkI9auEnoCGs+rdRVsItK+w+d4Vp1edDxY1eEgE8WGYajzyuWpYor
KQ+mauV6MUAOXFO4JOEakFYs4mhIWyjJ3pEU9Vi/moqIn88Oqih+LDadSBP0TzQlAOFSiw+FPyb3
5/z8hNZ3Eo4/BMmgJOpTMRjozNX/DPWnPT/15/X6B+nK2hlwyf1MndMHAlkXvLNca4WH7X4pmEb1
xtQ/FeFP7oSdJMs28Q82XxSGPWSXw7muH1XKLkTsrJ60YP5yTtCzZqTcJ/16nRFHtGx7IuzyL8gW
6bXQm1nUJ51liJcWACep4KYqDYMf4Olu0+qCmo7qAXXlnVhYKasKFFkoXcG+WB9vAj48VtYqch7K
MSqL+aI8vqC4f88FdaFWgvSgbvVyEkZCd50mxTglX6kd/UneTacA4iKEJ53Mm/7CdVsqKaEjHcGH
bj+wsWImYdN0CdvtUx5hT61J1rH7opVAu5VEVvTm99Cv1kNSR7/UTVRPES3xSDMBxq0Wg0R8/3ew
QLslbTh1LPks+m2NqkPEsjlOfrElOSK+v+dGnUT1rqxyFt3ZxLpPvK5SVBU6F/Lg35+BuVSufkJD
fZJPFEQj1tVIYZKPazI8Ne3ee5KZs/jhNyEdxWsAhBlcnYPAIrzRpQ1wM1QqQ6UZFA6C5CEpmIcQ
xoHW9MguZ5b445E4bT7ecEWFyCwXjRNQD1unAYJw9u9a9DLSatnpVUgDQOV4SRPZrFGohV8cnee2
gd/eWF5y/prBG1sTJ3PePR4DnUOMWBsQ54ffpvLG9NpL+J4xVHtlVFvIItRELhI8AXva+mrR1c0N
UxRInDzt7bgfNjxJLEoOD32rdSWfFvdjRzBkF/v8+kUoolVQDD67pjTEChfT/Wl9ZyCk78dWuNjY
P1YChNki2deeHw8bnb6YvaB57C/gXS1qPtuUdKZTBg2AJ8XHs2ZXZHGY/UXQqH3YHXqLTO9G+RBe
KP8eGLrVL53CZNnpqGGEp7yyJr2Xy8svXp3j+OiTQRxs9vrFjIbEUdVlwuYiLRc5G+64vkk/eWtD
eO0DlaMLu4X2jLnbFX0P4fGEnfF/2AFXLQvk1Adk1/GjvsShhpJIKVzGgETvh8C13Zdvx0EXsi0x
03mp7V8C6nerMCBOCoUyY6O1dNRZlPp/mIhOMFO8ItozLS1yChk5YiAWWvgutA54z71HKcuzwgEH
zIgM3D18OacwGn+C7YphZWixCdE0hrQtWLpq2ttfdeWCSAn24mhgZIAFLuVO9wtCI09b9LU1zIJA
6bWSGIE1V6YjlfNbLiQDNtSaMUz2EA6IKhaE69U0X0+jKQt13UISCqym3MAPklbkc9EnYGcqVYOO
pHaitBfnK0yl6axO8gcdw2UsXSI0MAjabHyhDne4vtHGOp0aNK12ES8O0JFTwIuqDO3sdgU8OMI2
LHRypbJc0uietkpEtmcHW4B5v9Mw09rfc/xxsvoDfihDuQkp9Era8EeYsP+nOPFw1V/STcPnnZTG
7eOpXstcDfFJdyluatcB6k8kNvWWPhw8xlT+StaZDMtTmeaHllHZMLCp6V5RBmSIUD6lS//k1ylC
ofnaTBR5fFBZGJQgYhp0im8+2fuDBDtrGkIpVhVMmuq+PJXDcKpow3zv2TbhEwLU4WpDCDhb15lr
92Bkn8vwDva3aNUmlK/C6Nwk2xSi3T6sQoQP/E1q+5zeTJKOXGsGXM+sO9N83mxIe03oo1ZtHOTX
pDsCm/6kUMgfeCzhfZdQ1mLzz3yasIhfJn5x00dosyf+BRB7ct8/KR+Hu/qA1mRnTB8YGeP9Bw01
aCvyMkK/3vWXxUcSah2TEwFqhvJhAK8HmCf7oIjlTSDHnV2h9QXqR+NN6VU3dwH57s5bCBg3qoAc
WpUMJHujj27pLSTFxMNArZYaFWxROMsoeHBhNf/KJe167XA8lGhTNi35Die6GGPvZKQ3NH8LzJKa
xzuodEZG6EVtqEDW37ZQYX9LZqQIqA6eRIRQ/UHMrdDStAn0tffCuR6rVJtdyXMiR92PT2nNELhp
0QrwQ3aB9QJ69/o1CYaQAZaZX+gAEy/+uXvAJq/8ji5amjudAnQtVhSpTIhIlQWhymbU/vy1PsLe
IPjnsbHgANWg+rru+4Gc8wi0NM337TkbXXMJqLNm8pCsLOXMpOjDXY8/EEzxXys8uDUsJZXJjjke
Y7nKO6VeQeEmMq2kEMGnKfu94OSdhJU3mYaUfCzqFZ3xO6bHUljPMjQ08PjASUq34KrDMVOrUaMs
YShQNiIXMrVLkMJ6MIb9woRqLPMvzCI1shp9hTZI0ZgenW/gCUqp6dIIKj+TAb33236+BMscptYt
2LbNwhgrpBcf8MFAevofAWYlfwJv9nuTmJCihpAQ71732jUJ1Y3J/kyH3MQj3Y5TUU3yK0+nF8ML
sPfxEUxUA6U2lZ2jjkOS+xfCC8vGkwqCpBeFrFgoGIre9qSZiRJYIm4iR6iOdK7dT0pOzb5p7yXZ
vlqeaGxL/gooZtC1Ko3nyf4v2dp7O4HZqBVI61oUSqX4a3JtMq41srNxDsMKl5Cc70QNAlqRGv/6
3nyrBr+8hAlOMfRQprgFmfDjyxEuxYpgZJAy2bZTJfgB3rpV/97GeK+x0/DTu/Kx/ZZYgOJbmpXy
3M3px5g/cRRT7UyRXYegtKAiqbyElOhT+Vk5QT+kuqK24HEkS8HI70nLkyXxSAtLbs1y60cAsGH8
0vilJekorDJ7YmIp2zOX0aJoQF02eE6rdOs/d/VjyEG8TCVtisrv66treMC3OLCONyk4MWfKsiCn
8ltJjymlZAA84MSBBEn5xaEAxHkO+VdRuunFyf7bnbVjKsKM86zQPNcIagO5eyVuvz7njOZby2ip
CPkhY5W0q4rPU+y4TsUJbdk17ob3yDtafRUBQBV/C8BPWfu5XQN6Jet1I5fLHYl7kTuNTbkvnXTE
itBpwBFwy4X60cOgZhcX9Q2ihUuypDigHaFQXdnKNfm2myQz01Lj7meo7FQih+6gGFFvHR1F/YLd
CgOg3rhwySBMSsanjK+850WVxuX8WRGFFxEHYntD46vQn/9haPspVA88V0UCIuQQz9meZBiTvR0z
7uclNKNlA2dO6beJ6QG+mgw/Ve87S6P0vBT6botzLqxEYiqfxPSVxax8OUbavb6tqiS60XHvZOwd
BtTnARIIG3QI+pPuB+gBpdRxA0IZs1JrUh2htR5Nk2ejVngVfXpredr7ajH+s2y2yfOukQQyXBvS
n12Opj4ltXpjncG1K10f5sTpC+Z1wMaqZn5ep0UAw6kAmns32g7g+viWp3/8kyzKRSkuB8dS1sxB
9sSLAJ5Otcar2BYuWR4P1wQzI6cgcpfCQevshRVxjL1x6RIDya9TPwGXWx96ZA09VG+FSVsafAUx
9THNIY6+GQpfivjNGQIZZhH2tx43GERwoFU61Ul82hNYmhRedzOkb4FPFqpoPM1i35mk+fDVjUGA
JmGYE6iKZv/kYKkQ9KMYoR4jUedc9XPkxarvIN1QJpSNsMTu1+X00uIsN3MWMqD6LXGGstvVRTvl
oZ0ZPlqzjZ/9EFJE8fULFXzjMnLbn56DrSNcyR/t+ir9sLdMy8rx6+qKANrhsKfkf9ISzYPfi/d2
K74kfPs7o2DdM4s5FmhnivkmQwjO48Nt4GEcnqZMzu+Uhj+4UMJ77o9UrUNJsJCYXwuWpHvVSC+P
WCtq50Qx05HzAmnq8rXjvHoUlPkzvwnUZ2UpD0DxBO1p3twow6BzpQMrYW26qCyPu9mNNT3YDnFF
9AeP2juW/4yIvqY7oIKyw158VULrAzEnvVOHVXuoCqb6Cw40yHaRFHrzYfk/73wl/MMrZBhlY9i6
e65nnqiI7KYbh7LDouXSA3zvjcpvjF8DzTNVMijv8+paboVL0EpkB1MjnDFkF+yfyANeewyCgP7U
E2ct+cnCsa7R4JgUMs1PyTfwlH9zmExOLzE2GIyQDr3yudm32cDYAFBVPdiHgjk+Th4ZUuGrOsb9
+EXDM0WvjesLyuZ/Q06xTkoJu4Ku+tDlUvspWXw24uv2fQxa0TFnANrAgzhBTg1rlBejl6NOLGmp
6ZyyF5I71Z51ND9DdlD7deDvX6V2KktBsv0RduR6XND0mVLNovX2euEIsB5loYkBs+a4kdChFu1M
Dlfva33ELu4+HDQ2JMRsAsOXhUQcZnDyCS953y+219DfLSanv4fLjDedRZ8FxEUW5WKYM5WJmM24
Cy+uahioKuyDDvPXhIfW46h1KTHuLJLPnVA1fL6bd65opEsfX55U/oR7jmdk6QRn3WhGNmsmy4GZ
5tJ+4XenxskNpLTj85vBpW/KdLHuwKwT6CqC6b4OiDzHx/7k+ge3f4eOzEWxqWSjb93MzanTncOy
vZCBym48gV92NP6jzzO7ijPzjRWCKP0iipkLekkW0rEfBwc4cCAZRF7cxOmcRJQ1nkJIAy5GhGhc
ySLAnJ2I/AcPN2LZyz6DxB2Q/9p+Z3MWIjr6Wa79PmaArWITpjC7lbpHAn80zdn30wqBmnWO4KwJ
0jjKvgzsQGoSDiPRdFb+00sNkwAwjznUftxZSVJyS/U3X/jU4A9nySnSYxW4GAbafW8fKENtMr2c
xX/vR1u+1A8XBCOphUzA3DBfXfzNImg3BB9rMQjKGCEapRvpSFHJtNaZD/nLVdkBrqCyDBDXtQL2
E/A6Dz4rJMbV8zyCIZnGTHUk5TFeeC+gVGxuSfIo2YXgvxiP8MMgphMte7Xv7NtLcSGrR7hlYrTk
otpQwJ8WAtZcPp5E/ag3Iz6+aZyzPLhS/1YkD+XC6qTnMAcg/Ed76YdVd3d+cLaQ83HThslzvnHd
sna11q9BF5mpXn2LPrt3iZcMWNwKvVz3a3WpkfAm8H818//wh+dxS8WOmYpqH4akEqtMoskvutEg
PdmOW5whlcfgoBNlKr97AzU3yEBzuznjvYX7bTTiXyh2mkUb+IR6qjmOhr6orwTtWqJblElX1S2G
WjK/RTtG9LveScwGypCVyykaiEd/dM5pOXFX1W4k/2iE+MjXn3i8kBMBPIohhrlkXCPPfRVbJJDx
XuC3qmx5y/GzP9NOnIuyJMIDr9VDd64y03YcrS8SB6q+h0E77d9fHrlydt2VcNJnW+J9SXNVRV2a
INpMzsDdBhS5c7f2xWiY2fGCjo7aYaLS2ZmEhf/130XsgaTCeuL8pVaa3ABdStLtkSrPoh9Y9Ndu
pKL8Oyggz1I+U3EssCpr5RRM1QpHWH49yrS2QeLA4FYQ20badAWFnenOYOXvPbznHf6m27uS6k0P
+f4EJ60dhaGK2OLvU3pBIxhamHIeZGWjtDyG4L0FAd6KCJwAdwHzz31G145nNIK9oziujs4qLTph
2l8qhyI9D1lbhx0BtJkOm2LSJqVoHaPp3NNRQVB6vEEkv+w6DZEFOPQdQTVL/8CHhZZ7/cka1Qyl
15KXmQfgYHMKHmzYv/jzV5fOEdI9w5yibsL7P+B0zt9OmEzc+7Wc1mo6v8aQ+mApKkLXD7c3I9ry
VeQ3oLc6MXKLw+BUw5J+WR7paW91HMkkjvChdgG1Lk3rJlDExI1PrjI9MyLkH7IMybiBTS9hxc6q
ELJp0h2RrCbrVlGIlPTTCayrJh4umseOa3jCkf7SmZUuOSLzBpuhNk1+4GVDmEL4dgi8TqlgWbHs
naxvSjXL6WLqa/a4QlN5jHOb/g27nEVJDrgDXHYL9mXC8uY/pdaQE9RPs7dVOrd8jwEMJhdHCNZM
6E0mGsPmJfmAvwS8KW4pAi+dt635vzY/1LDxdYdHETripYzuzZZkgPWomn+fg7a5kMj5IWY4U624
1wgNnXBA68xHcY7w5i4NEDSAixRgvUiPJmkXiidQNynhqnsA5xM2lTPa+Z0B7ytSOVjuDe+D9mOg
2BAQdAqFKt34OlN+YznIYYuYJaKgqj9IRXhEGLc9K7xQrRw90lZzVA3FLLCMokvyVp/eaBAXkJgO
0RcDvP575LGhiHB8IMK36nM8jYH+gWKV+HSqFy52mNddUUdckStrBs7SmDScV85gPlVpdXAGL0bg
NnSdVLPxlSQ2iICb2l8CgMr8dHc62Ext0XLOiti3q69CZ/2aOGbXf5GVeb8XnhcHgNxApqcEAjN6
rxcJUOMWeSeb0/qiLcENy4puA2VKxmTwXgA0PLlqfwJz3uVxQxcOlGVIssuIy5PE+H7flgltcKv2
5/xSyQf7RkFKJL5rWWTjPM6+X2phr2T+ki3EK2bmB1uLzoOuWLxeZy7RIhkPksyL16vMj9HunIJu
MVlzqCsc18l1/nX19ybf8uxJjE0eYu+nDrzx745JFSjwhxEhO6OEBjKZOjSsqVXg333rhO28Dgle
ZePNI8AWwGWnvqvqQkauzJhwacbEsrK+4TK3ZlmX17cXx9MnL0YCzpB+oNiD695h/aXECiGGpiAW
0PwK5xAdXFaO2ULWeRiJe/MI5H2o7Il9yBgUWnxMIdfuqOv0jn92PXPY/bqJ9ODSyyo4vf/3xPI1
ZniIX9RxsQVSKQOyRZziFN0+FZ8Hq9Sf+sKlmTKFnFvti1GD45LYPHuR2Nqb70fxtFJ5zb/Ka9bX
SIiEMFpa+qZY5aF4+HEZOqTEWIQ9Yf9DMcWnpySA5BSOqkAYXEfamAAN8SHGqKp3qjtL8dj4FCzA
KXKFpFcNHeu96elezHWK3pQsOe0gZ2DZ+1RU8OBidAyggDkRgcF12sZWX0O3r7RX9q8P0Xgh1hb+
1Rh+YqKERDBJQAxmhez6V58HVmoHbnNZDl78wUA1dW32p0KeSt3kbdQ6QBVYKFeYgBGsYdU7dcg8
JxrIH2zsB9Tj4MwgvorD0csXH3a1m9yGAAukUMvl2dZyrYg5xlgDKH8Rhe1+qaWMocB6YMQWYpiK
7Vd58xu8PlE9qYy+JPAdIq2vqlcUAj7C6lQhd1TRzeOirv/YEoJVP2Ych8C68WT8oGYV6zhbRwEX
ZRO37SIl87ZQno+s0uIJhyY7tFirbtDWqGD40JBry0lqhh6Ef4UFIqc81B2zcMVihVC14lnAs6FC
P1JBb/IHoe2EkDU16pvxlBhXBkxc7zMDYd3Ud7jgVFi3PREWn1dwx75GGvH72VsOhVY63d1C6zAn
ljVhk4WgEAEzEwYhlmNoS1sfDr06b2IUWfATnLTCNweBifqDOAOcffTyoLsXmGKSjrClH9ttZWKA
jjSPqJB1R9dhd1UKgf3jKwLYQvbJ0DQh7RcqH7gWnctp9e9X0zf45mxyWMLvxUTKsFp/7BKLDD37
tST7QTKQzq4n0i6eFhR+1aNCFKpkwo6Jv0xJheT9+rTlNbi1xSJQ/qMMoHpexYGw1tv1rUmo9WuH
aDh/FdLKHFoR16vYNhsoxO36/oXoSH4Ry7H0WzexNedWt+jmwqb3TvCb/6avP672OhrUvrjtCAmq
4gKAQryh2sGC96wTBYUB6g8HMED3vYiOA6SVv+GRlpNyT893pq0EaE/c16GvUZL7A0VsP4cxOQWC
4EMBK3RqXtRXT/vDCtRZrF+8Vf9HVkMzVySXR128AiUsi2yZUccKDSLIlZXeWTb6YlocRKvdFqL5
bYhjynHqrNrlHVMWzJOmwKiQ1gY6qstFiGgnjGyAkc+QK2go0Lm0TETE2Cpw4eVhBSrGt4ODO4pM
oo3gWZOAh+vx5Vy/L9Nb9tM/mO6WCvRej7/IRmHdG/6U4xCic/KZCZdavmplOBVmiXO8WR6OG1Q0
rTGmBYeeRT09s4d6RrMfMdfr4J/+jmsfPhWMdt7UmnN3LSBrlD6nwgZhoAQo1QMIlDoE0mgEyIy9
B8QXIGSEKnNZmCq6M3PGIElcpZQKnnN2Qcj4vn/hMZ7tg80c+COGosUTNfUJkaybOOUS3/Jn8Idh
cGZybzV9er2KbYzN6eejXPno8s4NJqhpaNwGy/KQuGiyIuLk46coPdwQdp8rAKt2rydzUDlMWNRH
fZPnaJfZZv3yn7PDz4KgiM5QJSs2N1ABE9Mvt3ffdQ4zZE4QtCLQzv6nS9lZh0MYaTfWE2yR8Oi5
9QzGj3lKodXJi4j/sI96cKPcFCY3N8/O+Cw5js+vo4fPvwZUy5KeMBe5W3uvdHi05hLD2ier31SJ
5Aqv+2kSL+jJMywDAbiDJhajCWZBVrG/tseVxMRWJvztaYWqWw98mwgrS2YxgyGNz7FnR1JUBwiZ
02/6FDHrxV9pgrFe2UKeW3nGCDF/ETz3yusFuowCaMBTE061OsEB7JB7Dkhku7JSEUvC+4fF6Ima
PXHI3tGhjIwnFROjzHMZNUEuTHwME6Z1IVcnO27hmjkAib6AWVHLbraum+2wkO2GFyFjc8bVghq5
e3rPMj76U7fFOuDCGH8uoXVD/Bfx6PE69g6ekMnYerKrZRj7psmIywevcqR6fz5pTSEPK0mHq1KQ
h7GjbDgWWbWDveo+NsW6vOmLEP27ERJLVvQkaEsmGzXfORYLoQY6R0cpsakpvFa+SpbvUXJdndxq
KQQo3o1+lM3PRYqCsk/5Wr+zovSbMVCyGPDrTzlW4bLKLHZYKP/x6gO5oudt0zIa6PD49d5t2Ybn
ZQw7FEtZx06Y4tI3arpvzz7E79BCLe55UTS5kuYTXnwWoezZ6igZt0K6wLMtEU9zPZXX5uSEltLd
jcbNeF5yOE29OUbURtmUoN4LArguYzSw/MPvIo1+u1Pkx+u3y9R3IS0hcCD0eVEny0oe77sV5rXI
EqFXUoFj6AHGMMBhzqOHhjlAP37/s4rh6P7RP7K5jAnfvxKXNCW2+8ghhWkrjZqkPO02Wu/NnVl/
ZHLYDPL4BoYR7bO3EEsg/4F7xefKYZA850ko047eqHVi8j+wpfw0XeqUUfo0OcE2yj415lFsXcnW
ka9v0SfhTBCEX4hiRoEPT+UOazDltd3XbNhXeprXZmg1DTR7jz+avG6M57aGZOQBWdcbOrO6NOQs
l5jUzx1KhrY95kgEQPqCt8BGNnSkhLmPRkYRFPWh/oOu6G0zfbZU+aEz4Ikv2m+tsjtuY/cxW85v
1hkp45hEgXcUPcshiF/jGkeuyVIVGQlU1nCl7NJKOwrYmklCqL8qo0FQQyZaEPQcycGvCwBJETXP
Q1YwEpTc/IPWgUuzOpSXUea6/ue8WPfMoJSIg3v24doca2Lqp2tJ6cQz4ZMiH3mFJQRTgDGonK0M
Rd5rhPlsVD0eYO76pz7UQ1rk7P+wcRF09EkP5R+qex72Jq/MgoifxbkwR1+iuvpGV+eDIJzg36xD
axgYfW0KdlSz6kB7bVazPhtTQ/miz5Pu307NDSp9/KlgSratVULz/FUI7jyF1/E2SC629FvkDm33
upyYyJO/Pvq0ISoK/lqzqK/kHyyNXSjSlcc90b6Jl7C0HQLRf04o+kKi8K1SaDqfBO96FWDFxDF/
nLwRTwsCCQhrvWL41aUHN4/6NLOUZfZEKkMVfTBZVhogNdBghOv+5XVvCedd7DjcDHjjXKnNv0G3
viIuDD8b3+7f7ygO4L/v2B7iUQ3WxldR0gYLVm3h/AZYpqG+9ayIJe+e4Q4VGHNmCrUZSM4Y0S05
iftTHqTT/raS9A1jXB0/vl8hW9dpI1xw54DxY3Ig+pUva5lzx8yDhl7cikC7VsvL4KvGbTAMqDA/
FfAm9YykYVF1S9lplKBY7yniwOhTBSYwhfPanQbvk0DwLcEHYdSZjwpjq/tb2hMYKz2WTxam7Jlj
slNFYjH51CZmtMJ83QLnX3wIr1Bii3GDNjBnL4ZcOSJpQb9W2XRBksyCNS7vaPxs+GtwKvOiOQNv
w4J6A/ggW49jC7hyfqAQb/vvGFXcdzzxVKTEx1FMrQi7PDLRpo273fhIKgYHRAf6rPta86kpm+Fp
+DM/9Cwk9iZLG321+TXslv9neDLXpkgJ3hEDw3nF0GBKAFAc0oSyzJpQa9RlX02DLsXvlaHpml8K
9JFYMFE+peiC/UZbSrcTVEEZY5i0UQmOWd6vzCz+Bb9Fgixe4Hz3z7Gcog8m8egZzDqM9UZ1cnTX
i+0jw60+RE4HKA/9ZvxCvkrD9GAf77KQrAPlEWTKJn8qLB66Hl5N6nPpAD2NwN/tKzGePwsdOVCp
Yteipq3Mub5fgMKBCrYrITy6De5NCzggcXacCy5qS79YtpyAyPEVe9HXBhB4EgswChR7F6gJUGSC
hHyL4U1NS/S5AIF3rYcNx3gdE/TPwexbxAB61Sf2iyPARdbdAfQLAnDtr1X8u3IobBXpRbrDbKVb
TmJgSY+4mdq/eiRT3cc+Tbbz/FXWcnpFlp4XyjqQK/VZfeG41GVR1Kt487nr1nM+yhUyDREfm3ff
yfFzmwAoG43OKG400RL11oGEuYonSjD9yqbRSOu/FgzWCCFCGJuorOXAfnEJcJH6CV9+PyIddnXc
xmq6mXPH05MNRunFsLQS88Yrpkfh1IF0whspOQsnuG0L12y4ko9HRMwO22Vec8WpPkhvAclz92yu
TfVhztTgFWA917tAN2YU3JfZZGk2bErAOagifJZxD8aOcPHJydSzSvp3MZasVqKCnVl/Yp52ClYU
ngU2RfaAVd6u0DJO/GV54VZzEhUP6OBobgyVNvgCtIumiKcAcEZFWt57nES7S/3ZUIXLZu7kipcU
rzOm1mYmeo9vsh1xSSqkUjK+jLq4jD9IuPQcwUH6AmHbGjTmFYm7CUbrKryUPyUHgs1nhgsTkdhQ
p2g1C1jskdBW7aPhmWJTW5GUV+A8RPMuBgyxtIYBl/3nKG6Xdf9yAQWYUBJjjAmpVRBdOPPR9o3I
cs5FF5UgWJ4+o+M6PazEoRwTbvs7YQb/GDv1oo0n1sJYBtWROhaj6PyVNBFyLvAu44J8QAJPf+Ye
sm2YOStKqo+YQ3/ESM0Ql511RfEEpMFtavTinh7IpnAjYpWcXXF6fmgTQsLB09YYCtHEDCH1xit3
tfN3z6H6RZxYzfAfJJsWo+Hd0n59sbDWIx1KuK94fegxDc9m5zMnwFZDvR/q/thuTc5fe0uzTNdJ
/H0bPvUi+LyyGDXoQT6viXzS84QEpRbuHHn3D0kyBC3K+wWyoy/ZEmsAWjSx92usec6Ldd6if5in
pfVEr+cJr7260lJYws+Ae4GRiwQ87yCVeBGvvA/GXfeJvtxer6p9sbcX8ZQ7NMfSXb/2WPFWbqdG
RXHHxlXVVP0ICPtBz/AEHHAazBK4k8gmE63Pc3W472pB/amFyLUJd7A61hE7trUGm1xrh5d85KKX
6NKQy3qT/T7PCfzRgjNULrDB5AjN+q8yL8pjKR4z4ePr+4xMXbhZGxqb5nnkWszMPp5r1wA2Xf1a
8phBT5ICLtHe7rpFRnOoy049TVjRFO+id2zLbm6omlhrfz/p5QsqSvZukpWvB7QvNbtA2YRjb0+H
8Q+9ksItIJU61HvyLsNi/IPwB82Afa5X1DaHYpKgnra7K0AFbpyJw0P03OKTbO0OqegyDrVqxyUD
bk7/C7dNXKmXGSjQc4TKbccgBIGk94XnqB+ilPNjWrmaCEYVPzeA4lyG/QirDCeOvIbw2kTzEg/X
c3OfTBWuukIbIKujWKiZPcS2uMG9xQo4jPbZBtR8mCxDie1wj2LG92h13jS/AtKaklH81bUlbVg+
0C9vYZ3z+gZQ507mlpJY1D8cOuIJlmcSQPiAwxsSeNMumMByIF8dXiiI/Wf0aeM9DzpWju8sE3RB
A/EvaGsD2TFa93+G6WSc7fCiMP900pQOUECtcxygxV7YHrVTVuH6ZpZwL6AJ18z+QkjiCnDuDsJP
5oCjHu6lH32TMxErblvvGmUrmyeQ3Z4bZD08xpPs5z3Gxo2J0fuc1FMHOJvgBfprJsRnD/II2AYe
vZFzshZiUUxrMXuRxW26GbY3hHCJMnlgQ0g98mBHBJGu/3zkJFeiU1Gi+c4Wjq2RV3AStMZaWHH7
4MnT9JR7oqeYDNIHfF8rlExhBUBhRXQEnUnJt/pgzJJ5DhA98UxoBFu2SJEAzoeItBhqL2asjqjp
tyoQbjs8D8T4VTbI3JG/p228XhZL7TduenO2IQSGS4KaK0F8nY/Hk8VZ/2AuUw6gZT7u+hwxpaT4
nYT7nyY75NeKd0k/nODRfqpxxedSFLM5IgAx+SLuKptT6QkYAVoAk1qiUay6WN7DxSIcW7xZkHrE
4dR1ozOFMVP4pltym3gV6r03fawMzxNLsTTcnZICXXO1hHoM7m0kVlYocJWlyL0gH57sdSpNoHxk
/TBGcwAPRPITT+WplCKmbvZdWaszR9D5LZpAtQwrDNNNwoBUtJGvYF5/YhzDH2+vIp0ikEsB44MC
6KtrL6L7mTvg5ggdPWzZ5h66NFuTdlerr6LJ1sD+MpalY6p+G183UfFAIdjqQaRa7UEuvNpzlb2k
dtu5zSOSrpH/Fknl9EtkHQGX69a2fcvheOXj+KZJP4hWhVW1TduaH/pYXBnK/o3Exgvx+BtvEpdF
tL/whhn4+iSJTTHLebqjsLI3Dl2dR3jUBk39q7HhMQwidyDXkAYq9nQUUNWcnE2pYp6hApKCyoga
YbeeSg4BnoK2qLqOK3QKQiHnTNvSzS0JruaHUN/2L/GyLiKXvos4zxSDurREFcFct9qSVnI23woy
ZTio4QzP/m+lMHNeUxyoORQA4vA4HQzmtBGMr5qhf9Iae+7btuaMQv55BkAS4XlvV026PjT0Ia2A
RvW1AvP+IO5UeBmGbjoXSilX8AFExvs4djMgKwFRxExMs48Dd2F+wUIFIx/sG8JupbCBoDA8jvTZ
HvTR0FREEdAdtoHMXBNzIYNHKhbetHJQ00YVB3aRSw9pJB7u7HOX9kxuoGhFIbkFw336Ug0PGiFW
sdapFVAOoKER1KgTO52RcL3YugU2sn1httMr4dXbV52G1smxYuWoamjx5asO0smIiaNH/0+611bi
9oJuvXZOXZaJ1q571J/iQ6fMfIyKjX99Dd4plJrda5wC5bmrKexi6hSm6AWVRlWnzwYOP3sMTJAf
wlHEDXQ16aoqI+NYobFZp8ALytPo7ueEY7a6zuUJ+i9Dcl2nnb1NqCicY+VU9p3MxP+vR1Fv1ELo
O+FvQdEfOGNAGk9X4dxtwrJVyJZbW3vp/hsF4tAq/eJsr82qRM/uEZNnZVdJYKDQ2XrapIvBcFR2
u6kLO4wyHIZnRDsYXqwd5v1JzGvzuMMMg+9kaWAH3SP9StOE0cvNwu7OAhnQe2MZzF9qmIEo2Jm7
DlBAVvuddDMrlhNLGVxh/Ti5xRF0PHzDWMiW1AZIRgpQBOXDgu+Jd66oT2bUUglAsL1yeN2q50gY
f6pWyRrBe+paK1/IRf6W5WX+3k6+4A++/80U1K8DvdRP6mZq9y5E4PonES5K61hoap0QWSVDUfIM
qP2Lex8AGMFdk0AQl25wtxEwn8ywIfRMK1EL6TMfxzC1RB7pRVDbbRmrhGIzLuHqnYom7JD/pjzz
8QAZNgqoREg5SOylJ20RvN+Or6uW7POyZ+YwT/RzVU8JE5ZGqlIWQm/WbLtUN+SecOOGQNg+qAUv
7waMAiD8wF4gsgstwn+05uWFSvOyvQ/c46etJF4mZvDdy0OTJX9gITxND6ghZS7UjdlEUZndmdTR
SWjCz6dNAdt4bNp/p6HspjACQVclsdgHHCLmq6Y9rzK2ckwmoQJWGKRdZDoPebM8SVDvfezUo8O+
8hKY6I+MJTAROgdQHAFCix5rroz21SJjzm6urnnKuP8nX7wbbr0f7l/sM6Nx0ezaw7LFw/grP11p
/zCWgzA3sWYSh47OwWI96fXh+RiRxOgsBGZz3unwNBsp20O1mQFW5X3XahUHGQSJY+zDrMHrNano
TbNVVwG/a/6sMGF1zi7Nag0jRBmGsZfyMpsaAK6aRO2SgrmxbIbWxyCMul9Q8FKEcghbsxQbon3c
Xd1cdzgt0Hwmqdua9FoyqaCwKeCPCou7zMGdZPCqNWB0NRWvPJGBmLgJ5bOF1CK6zOeSxokMAN5w
Jyho7teY6l4MVBQ/j4hUg1FluvAhZUaiFqxw7Ga9LbeU7JGmb+3Y6AI797UMA2Id6aLU8anP4ZCU
kz1ZjORCxVqS5L15DpLFHCIDfLSffQCb4Div6Ps5XFDaMWJFfsfFBoeIcp2wbW2p2dgZ/G2aA0zJ
7iJwhAAC8J3Eu+YlYikI2bXyqkPu9npXMDXHhQGsJXzFDdK0yB5OhBX4SCpFc0RwDzmjztAr7Ult
jObfEK2g9K75oxOEGmorSwH2JOjpdM+BoHin4LYSRBjtsUi5bcatjyfshLaQAd3Zb3M1rMtnPSFM
wP+w+9AQmRB3+AKYL/S3OLMuBDquqpQYDzZZo0sWLxhqmda8Pu/MF9tLQVLErZrOxCg7EEqLORqS
qGyIjmOlY99o1F7pWs6W+8C4QvxvdBHxIZisTrwdcqyGeTNKIfgEoIB5sZGbshBWxN9Md1Svh/BT
2Y4TfT4C6ziwCD/qELZQtIC23zIQN1j5115AQn85PiRTIItDL+peVP7pyiz1dhTdTjarZWioJbcE
71uuzyuH/ODtapYxil1jwuZg0FB1cQD8wEQ5wlVPra7JGZLkPCvWYexdNum/DkF3/T4RBEjoGmjd
ikx3C4eCt0E6a+fzishbul71IcE9FoaCUmQW5NMNg5jZvZuEg91rZawQQT+QfkL1mwfcEaZqOu4v
vC79ZVk9wcxoHavslgyku5vrZm2MTaZUShkLWk3KUp8RWtPBdfrcSh84Mx7/Q42601bl1olFTgDF
N1luNlT2rUifUVD7IwK+JmCgFsDwCURJNpuGxSbk5Ctqx4KZH4CR6S/kG+WyFqKxzkIYolY/rgUf
H05y7PjlY0BT76QWnkggSImhzXFnq1+GiuQmuNXcd4BucfcsZnNzB6pzWsGiwk3YE8W4Ja2wTM6w
Q3JTTdoeI7UZ5FHEK4OmqJQ1/Hqa7eA2yea7L1divSpmAEeY7w4N8+f47itMCaaX9dn27LtuF+WF
U3PM3bdRQjkQDJ6RDualsZ3ibv8LmR6O1gBzzb4biPagYrH11L69ijFD7u4Fg7Mb9qptmXktb5tw
rBLnRFT3No0/XfNKyv6KPDPDzPt1Gl7M5XF50R1TH1B12UC0WMFPLqDwe8ifieNKMM+61t+4Tclh
Iix2BjGLg3+VOKmTefvLyPW0mDYlBIH+4YrewXaJBczTGcqjDlp+gjgyMjTkTadOGFkN+PxQElUn
8vC3I+Ir0lv4CFtIRuYzHZxDYz0jRw3jWHEEKZZTSlmNYPbpQpweXdb0bYlXY1I1tdpXiZh+1Rcb
7BZYWc7+x+mWUVmv4e1RNkWxxvo3eA6PfL+OTsxH8l1/7LXAdrkCi+CuGCpBZB8EJW881sgPZhaT
ElnCEvx+HxKtMhwUvFKSS3FtiIfAK37qtRjcsdoZDeoeiRiKEuJ9DmvT5/7HPcUvsRJ5KTk/n7QU
dNTNhfqnMDqs2gHTEkqF6gSTQ9yTFA8gx/8TI9ghH9PR96AOZMSsxaK9VEZoWexG5QBBNMjRFo3H
/fmsV59x7lwdVUPjgEEv7S3oeV7g8lzNl8HEa/Z+gi1NjWdWsCsRUOuvNiFjOEZUwY7oCA8bu7EH
UjShbpoNbOg62CwJYHPwPdHYHNfMNI8CsXW0yXa//pUJyu+uDG3FZQVuCQbE5EsErVYKhtIxpaoT
v02xIKkzBQrhURhDCsqiEUKjmMRm8xPGDgyUVTHnMZ6KMEi3zUqsV8W/B8Kpmgq+MGDniV2vIcej
bXPIJFNxGKXSum5HPrW3dueWS6z0MKC/99GLk/E6xyoMwNh0r1m1FGioWtT0uJBKPeXpT4q3TSB9
as5+/vmmt3lbTG3f/+mBDVWJBuW3+2XiE9Tg+CMp5sCcoODCF1mm8LLeOon5I/yx1rq/oK5aV409
O90GTPlpgJFV7m8I9tNXBT/lWEDoI2ej8npMoHGQDCoDO4nhsOURtzhjE/fcRNw95Kt0auQlUI6U
bZNZJDzSysGJFCcL/MTMNIQP+tOyr+y7MvqzpP6RE8t0a0BDv+/xkCfl/KQUKO3XeISB5Swsq6/K
z888DoGZyJSVNsFp7NjfBa/0bclZqgpI6vMHhe186LXnex4WnxGJ7gYxTDJwHRLIFc7FojLVdp17
lVBStVx9jrKhcrp4YuCY7YeZpWsIYMODT9OdEQ5kxvENnE6bdxckezKfbbbhv92aNKwI9pQzP4r2
hZ6P3iGJAoGPpDpu/02bLPAVmXpqO5jBU+YmE/zlMyVcEJc3HToBeQXebozvvzbtfTNtaspYxMT8
ZIEGXaZYS+/sZNF7PFwjreNlgDj5sRiP/LCHTEpgkIHWrzSR3/j2X5Ec+mjlhJolG8GQkeSZO5IC
0UbN9XNOPpQbWmDz/Qg5GtX6PYcTEugbExPopGEZw/ssBNQrMnUjLuxUhlL8KKkQ8e6Y4Re4f7uA
5ZAO06/2gDjj5bG+L06bxUgkld3FahRO3Qk7h/qi8j3tT4R/27IONywnraTZpRuE+dOAtkpay8vB
WfeXJCzC/hE422QAWDXOM2EeZZo54r0hvaAL8AbiHQaW2Aw/nTwdciBrSMi0VWMl6INTsNBl+uwj
iPMuol3dpliRe04gIh62Vi4hxVFQiex1H6PM9S4A7n2gc70eLq6a+aFNL0+H29bkA4Kn/u4uzKM/
DxdqNGHU87u5pxbhvkG3gE3gljFwQR1k1p0XanFvxEShqv3MGp6PCL3nR67Pc5nL6BG0RQkXmUcD
2kM23GGqv6WzAGFdKGMaMH3Lv7D+2ogkipk372KEZd0Y4Eq7ncp5az/yVZwMpRBlRhscCwPEoq63
Nc0M+lbs0TeAKM/qP643y84wqNGpIXO2Vwy5JE1FhUa+PO/A6V/YI3shM/QGmcYtyAbCxWKYr7tA
sqzTtN3vErLu8O4TsTc2e7wTBfmgnGZNdAyH33cJatTrr9IfJ4jZJwhQP1macTOhOHo0MOcsEGtH
N6Jjc+blZduZYBibkb3GJhatJ5tziBUG4CPzd8K2dFAaYlYVHFs6gB6krX1OwCycGQTYq5yV5TvI
QbwNb7zmCHE+ykxmNZQs5ULBvDAFsq1q9+tXodv5/q/N1HRQfW9XtmA9bDZAMa0AByH+jb66wDkH
kHLJ0MhlG9gvM00EP2oAJZg2r9gDVgTKOEYSLUYR4q3eu9tz6XQyHIlCgGXkheHJxWCXY6GOKfQt
E/OoVzEh9LicNEwNUw9szoqSbVS4d3xK5SWE+9ZIJHJTiiishWnQAlGYMGuSm/EVywdSYPWxkegu
11TEHMWq61CbNv3hYp60ONggueLVf+3IlwC941C8A5pbnb+mZY8YTRFV4ubEkk+Llo2LaFGhc8Fr
psOmQfztiOW+yGbv8CEQRaIYfxDKZZW0XV1Y2KfaJXkXoPFKZIPDch4iU/t/b0zKcVYsX/ug2G0V
u9flg/sKQAAXjA+epoDr2a2JsRgsuO+8CfyefcY1r3d+SC+TpRPrWbb1swjnqVKe1sNpMuKRb4k1
H577PZhNuualmwu90CBIpNc8h+bf5eyBysToSJN2X3cn8U0dDc56jcr2TsvEfTDFWq6QBZ4xgIxf
He/02wiiRoMD0x5xDgS8IKu80kWmtsKCc9ooIFpS7D9ZrDpVfAxdgUTlczz4VPelcKJebZNUSkCg
2kNAidq7vVCkLJpVMIXiTuAO16iN2HGM5Yp/2wITZb0Raz/sE+r0US+0ZnGaNBgsXwOOPozxrf5l
1DkrDEnH4aetkdT2vcSO/G/Q2isDx9dHx55W5PVByrfOzw2TSPQpBqMyFm7iSz6U7eI+m+iW1HZ8
gvIh5KssJpCT3RmeG4zB+MlsWU8xIoa5WnG+5cJWdXTr8JitAmUTR6TTKCABRFh6gbJzixj0oPyQ
rxfSLVQ3JDMPGa5PTkV+MsqNkvUpKFbfktmZ9Y2WGX32DJu1glo/DCWAcbsp5ym+5RFXLZyU7aX/
wt3jN4E6Wmq57hYQQCVjBwYaJBSdzvoGVUWlkrvREbDeyhXi1HdlCLVDoAAnFIOQNNeMwWWOFjge
ist6eDcEbOz2/wMFfFiWBsFh6cMlt/B0dNLHqkObVubPLgkAvRBm17RfxSlzj//GfVZPvKy/W8ZA
Fp5Xm6IF5pTuED43zAnbqmhR8A7h9vKVep08pVXblSXcPr9DrpAF/VeghRgptjwHTKGHScpghXr+
SGRmsF/3GMSG5GwXp9B/2qFmIH5HxbxTTBjx0T6kO7ILFl/U0tSlrEb4b/gMOQNKJJ+PRSrvwUaG
fcLGuPQsEH0eEPbrp3LS5fojDYjzdS2ZPzaoPCNE6kAHhmD7vIGg1wnhufItB8vmumhOBlhnyeGO
RGV9rSaNqkGWW9uBUkLWE91ifOuZ0QnVDURco5sHDrYB4pLhqsNjnDQnL+OibTIB/bsO+Rvadovs
0D/CNajSd1X48E9RVxbC3nJp+ugKYbZb2mM4NH5eFbV3wfsTh+Tktdnrqa/6lproOoniCuoj2iZg
QoEqad3k/KeZnFuLPJFmSotDDXbK17CzXOitGSeIVTh17xoTBcF8Klt6x6pbxGQqLkmwE6YoGZHs
ikfQsgIpxqOduLYOCRE6/zkJToErWTyZsAyE/B9w7+nJRBA6HGYmL3SpBKT2eivvJJ6tP13ET6ZL
Yddbz6TNdgrFupvuFR6MpX0S+Uq27Vdx9euQmIYQfqidUzxZ0ezZc4spz6tf8u6SYljV5ovWLsfT
r/DrxAKIAkJHbsgt/+SZa1i9hB/uWri/fg6WFzg/M0oP1IodoCdjAFE14nxJzWLGpLhvwYedi69g
8M+c6OSp1taR7MVTTvecG3kn3A0XNGlGAxo+Iz7yQEBKilfMe3lr50+be5sfxDUZZitkIJQ1t6Gp
Whzvt4IkbD6gsZBf9cdWH/30TiuDL5z4Y+YqsAEcWEYAgoOp/BPJStGw4Kw8nNdQc0rVfuLlBxkU
+clH/st5ouf8kZbBfNogt3xhsQWdPsj4msosy2xAitvNc172UcLqtbhH5MHrBgg+xQIJvxz6wV0Y
wIfmu/P3YweSaW4ZBYZNY87eInEbku1csKU6AIIt47Eosp+72o9dsW6GfjKiIAAI0SBvH2bsQo8M
lJjw3hrfJaUWgJ46S8kvL8ND/DVXjMDxj0c1cAQBWgg1HXOg5E+iEVQ/tQ7sf6kM1i9E+Az9WCHQ
ZwEJCLZvdpmx+G0iqShSGt2hV+2hAg9jag4gfdde8ALrEGzg0QrDaini5sU1OvNkPA+WQWYUxv9x
0dlU7JjokgLL6vMeP69quxGFiqy2VmNIA4Qj1PeMv1Z2nrPTW7szLCQZzgdMuDYd+JANjuyqhn3V
conYtr2bv95uRtjcDBAGasvKgDwfAaoK6tyNhzulGlq7u3Qvtr0fBrexl0auC6A6pHdZ3czomGxG
Fe0Av/bK7La1XZevQ4Z6Zbpse0dSp98UiM8qgmirtY11ZKxWVUj736C04TcxUYHqbALNUrbGrjKj
TknD3wxka7Cn7sYb4BJ1KgQ8H3pfR0APnHwXKYY2r0si0zyN8/CV/BqGH85sy97blONlJm9hpArm
eI7xcyG+4NZLq0wo2SN4MevSSkzqHyKmsVUJxhxO4M82di6nQgE12WZXdaZLnCYMOKbAFqPa7T8a
dye9qjipa0yzJ4PfkfzB02hiABGwWQKgqNvSEHq1QrnmZATYjJOFsyP1rcvveMMe4D/g7dZ29Sfb
ms0jKUNbYy3q8k+Z/85iHkwk8g6z19t3o3fLWzcuBSJ5l5cCfQvSEo8KryPbNJ2a8a7GGLGZTx8X
6JTGUU0XWfCmmaDv424UxS0DIMIw9elU5xHoKAVtnxz6M2LlK6bVpOCkfGwxF4a7e5j40Vy94Lyx
D65u4Hbb5J5wu0kGFI1ipggA362ZHtAKkvN8xFVC32ZFfRIIbgzrPAU0eSh5Am3CudmVHoKOog7X
nNOMJ6ScEphJUMfjaGqNsM4AqmfDsxCiCd714ew7YohLUyNeZNGVrPVRnxGW5PN8IiSwNOLyi8fV
yoosBJCwh7lxCUtzGO6fe/NYQvktcdDPUCaEoOELuJjQAKs5vmkqLhbR3wGAp8DGUYEVKSSWVMI4
lG7HlJ59tpnEzVMfe6AXExzJGTRR4IdzoVBoEgRNlDaaxubPLMNet7P8fJO4WT1ECUkQ6fINdXhK
uECim89q457AL/YGKOhyOzXdgWldGgbvQoSWAww5gOTD7jjMxRYps9tHXHcsZ+NlTDZGSmp+TkjT
LMkeL3OYNJU8Wf8oyFmDy30HUkksYtxcLq7wOL347hFsIo4BITWdIoO0+dPqD4OH6IjgxKx96HFV
Af6OYbKy4uDpYa0/c2eCGJ2FRYleJWamUr7ynVI7j8Q57od06c6p4KnZv0JARq7CNXXiAUgKRKhl
93/BsqJ1OKVnmX/L64gIr5rAgrYFf27ZLEDOnow+MBWDTgdr5vf+yO6XKicI93twiPAvPYXlDV/B
sLA2sHOOluJpz2TiwNXYUQEiKQWDrDVDwupUIKKPkV6MbHD6JGuYvyxykctKv0HJos5fQ/Ya/GrK
0TqHAvPiteLyrGW/SvOWM4dTTNJbYvhJ7mwxloWBFFvuleREg5StqtRMgkgPcp2l+LFlnzCsKm+2
yBz5EATu2uF7HGXjPu6eEiv5GBXqUMrTzrbRRf2M809hrnkI16wfXXG5+1YU9jD6Xx/tTS/K/hDn
IZ2vCDSg6+eAfoR/90enE05dcbN4VPxL/WvDFkuWZtG9j53TL4HOdLF2u6dp46AbhEkbjKwHqs+i
+vDKiYatCzHu6At2X0nyVDloOXwKRtnAWOpOOdSS4I4dwoMosoQSqwX+/MxSd3BdC5K+dw68q1Ry
1Su4v1TcL7GhovuoFPQV0ZWwLEvPgbDikAQW4WGojavuMjZRnv54o95ZV/wQ3FEFjmU7zdZn6X0L
CormvdH/vYTjSEYAqLhZUz/SGlH1Yv1aRNy7h4yJZthaLj89DJZ0n5nVF5q8W9q5eYlzBlJ5Dohk
sR+QXOYTrl11zp8Qvq4PrS88riNsRhEB0blaWMrCZ2CHuFz+lMsXpPGHwX99Ub6Sa/8do12d8bdx
sICXbC5sv3V0xpdTCT5WL7J9BauY+JQLpw0Zpc7mXIhrrdN8QGZNZAgBmj+LnnE22H4G5BXDVTr7
qSPNnDaPZx8jv3NSWipNxJTDxGKKflMilfOgaqQFvnZqnByAZ6AK/SEITliwiCS9ajWRFBV7bHaI
iYS3mOGsJanIwuHGAUUldXHQWFBQxmGQv+ChgvJnZfpmnItMBwgVsWHO7bzQVgA8kqYlI9Sr9+TC
MN4u7h4NC/7BSK/hiHAmr1KTBPP0OUqnOEHqomNklkj8vJTcCWeiTzTq9t41rf/ELwA++CX4PsUs
haMADjRnbPzy/H4tW8qZJNBF54z3q5TmknfQdzrTIF71kamqg0EANQiUlQTUGZA0Yb3EXzV3L8NI
cOJO48rz6jUFrigxodzsl7pIQh/2zEwFnislUgYtHd+HLcj348+VCiCyFNhD3qI5RY64PAFwwCVK
ET7oNP3AF+z63hEKJNssR/qqOkcvk9/syuDWg6mjJaHpOtqqtOiNAxx20NK9AS9Lf40RHV2jEjxJ
olbJ/U2sQc3Ai8U+zmv/Zb9Td81XZ+rjI04cbTdKG0OtR6P1IMaw/klDFbqLtMtOdoHaPjh//k0q
xOH9GeGBK46yNFB5NjAzOKXaXts9MQdKQ4FaZRrgc0cTZNhdz5PX4sdw96Lfv52x4+OGZzXMpMbT
yIePnrGAi0kwxBYJ/MVQf3rIpR/DIf8pFbDVCI+GP/nRW+9p6+afZxR9DUsFkj3+ViSfulWjp4oM
XPImPmlyS9DYre8Q8z87DiLzPp29K3zTav/fq5UVDjbzJOMMW3Hzsu6Hw67k7Cmce/NCLV7YYVc4
bGHyHZkytGbGFnkutWZcb5cC0NkMWvGKQ5sjr14bx6JmLxkR/siyVp7Rdm2SS+vBS3gX7hDlhbtD
+1lUhh9JcdzBvCKBpzxDI/Ri/HyJppJI/AaB/rLeNb6RD39zZnd+QGOO+TI2UYga14dvPKtIntWE
a/JYkaQI0lkopWKrngWNmTda4AZ6gdrPqz2Ce35QGd/oOb2Mb0J18I7f2/X/PJyDlQbhaiUh+aV4
kj597ml9W1EjRqeeKE1QrFytGFCgKL4vND+wJVNRD8tcSgakmKP+RDjeH7g49kSJiTkNhWOk//Yh
eC6CNM+LP+chW+g9dKYrzZ68y9QGNZaxtLSuFflyXXBcG2IBnmdHZ28jf775LBXZ+PDqFVTAUc0g
6PlgLTGziTz3Q6XQzDBfXnuV8vWDCBecaq7vmpx6BpB8jLA4ELaIIJjlbJS4CKc2hiLk1222xXQS
j0LQ8NNjZVVYkII/EogfRCVsOZcruJWfOnhOI3YXAJyA04yfIqg3NTyOIhAYKOuOln0+MPMR8Y7q
+wHqGYchpJwc55j59fOlVB1BxVYLvtb3m4j1Ia+uGE3u4tYN15hBJf7OCddkOh5+bMl9ahdVnnrW
qsxXYX3rhz6LoEZqopgDHFwtzbAkDSjHzNOmlh3nO+KFoVb3+39x48xZbtyFq6mSxNgW+arpFNmj
dDG7Ks8kVLBb463FuK+ulWyaMFafx6a2nzbNaJfV+yFNkYGG0svWSDrUmy/5QPQHhL8y0yMilSSc
PxUIhR8Ihsw2oVwcVixcLpcEYcn4OLDAoMQ9Znqv3DcbnwsjTXQQRGCT7aizWIL/xV58Lnxdutoe
yh5Xq+mgP06eQHrx4fN07DGMgQzZMmawskXtEJCSsX/PQSpF6JiEf1qjeM0CqKCt1efh40AYRp2o
iymnwl6tYt3rx/Ezx8DyhkAhSHq3i11WIHoS8mm/VJZpAuU6I/VFl26wBJNyJIRcGt3fGMbzPD28
0kwacMGmOyzooF/LTOltiqiHgO42mNQSLHn4jKr5lWn3A3L96e1h16CvYjsyR+/3YS4H6E6JDDTO
tMp8oXJyAFhGBwiwGGeFDNOt/ztDXbVepeU8WXPJxPljoTnovF7jBxcJH/bWaNmDcL691Upxb0Ik
ZwDFUOCCpvokyrHgaPFj1XlZN6EGUTiy8TybW82PlX8f/6KbJ9MIrqS2eMCPY4SfpFQ12IdMUnWL
TkJre7+8GYd7Xh3801Nf8TYuYaD6UVgXS3J1kF1NoPKPPAf6bBzMCI6kCTuiMDLNTf/TNMCxivXt
s9/rceZNGnBVMozHUo0CpPa44QA3Vw1UQHXUoNzbC5k0UzIGCVp88JRjmys516U0ZIOzVVwVhr1m
W2bW0IJQwx1Qy92AeV+Is6emRxRj3FQackP61M2Z2OhVa4aDDqBRo76oBvRZSKFwh+gyvErAOsSr
9n1hJA0hLuYRuKez46HVxJJn/KBKeCuikhfTnvLdNUb9jwx97b0PA+yPrKnJyA55GUsXjJze/uMj
gvDvMCl0uqNYgHYRbMvWFZZebLhkpk64cOKb4mY5E9B++b7VPcN5NI1FKmavgoIMZidNg52yOyf9
m2LZKzItguGUDeYUMLhIPbSfLXtNiPCdFUJBYDnJrTt95MBNx3XL3rAdzI4SUZtfZe8qPxBjpWjX
0rzUPMetFXz1SHBQzupMV6rT9yQpL+d39dQ16h52fk6FQcmUe+uGQyglT9C2i+v3ttzlWTxqedxS
p+k/5fMLaJCXub3uXzJqArSfSXjINtZPRYJGC8vQESIaue3vnQaw556bWyb4L9oK5cI9y6munsjj
2xUrEnzDAEypgFzC2f///RNT6W96ycAjWFm58MnCYofbhs7zpHnwm5IW5nXzT9p598Us4e4fKPws
mxT8lrje6eK9pz2CfeK324m+5KGrF6JLsM4SzsaNG0WMUdWM+wfOvxKp+mctoew0AFHBYI4gEpxH
fVHh/9YJLY8M0Yxq6PU7o0/UumN54EqfM0RwVK4xzOcW25hJTYddNXZC7heMOoV83EOG2OpeWhbA
eFc5vzMZxhC/WRlaPUMdGytEk+DKuOcDdOO1HZWq3T/0uNMTgpIq/VeiQH9Uq/wPFDCgqJUabyPE
3uzgS7Fs6kCYNdbGiFIPIZTdpqF/wRkdLN7LsdCzvw1GkdvjyHG96bxPJ/IF91YybuEOAgJ2nULw
B+a8pKkS2IvMDgGn7u4OqZaMcY7sG3lvqzEeeeWPt9qwIaeH6JVTbSwaSwSfxEBiymRcxhIn6BfC
SzuS8jUhJc0di9cSNYbUYJp9HtwZpkUs+DNxqbWb/oYGGVLpQjJgbt6iywWXmuNhm9nhCjLl8+t/
mJAhSmnPkR2oPyPqFHly2Nv6PcnPlgdaaKImPqFHEl3W6Te/YpHtY2Nt0/4AYn5Zf5oE40DbVRiZ
f2iqyoybfsCvVf+qecw7yUgVCLK3yyGPxpbHZXLmflhP7wMfU7BLD+qvDi64IV0mVIhy8cjryX7i
wbwAprJL5jg5kCUP9pHd6CxgSqGJyxkpEyCvjNE6J/2DqGrso+dnN+bHdhrFkyRJWnI3CbaTca3f
lCbV2YSsFuLo2PnyOImjacred+MRbgAsXRS6vlgYk7KjuZ0zyg19n83uGpLByOsC9yV/4XwYZ6JY
p1oTLbYXkDW5aIlwOSiCGlFYIBrkkA9FOF2RhiRmM0V6UnmIKFXwjRL2PXzbudPCwVVUg9l0+Hfi
2pjr+ecpu2TY73gNWfz6JYdhjyyEEvQaUkNYCPMXYa9aFwlFA077I2egOTBXADgNLmXtFEOQ9z9y
SMvjfvRgGcevBJyRH0TQ9sRoxW7cZhkHW8XQ032gYVKqEoKR3kS4x/JL0OOcKLw5BBvomgzYshmI
gkpD5V2ZIzDwx0ZN2keGDnBO9Rx4QBziKxxYTaRoiLiaw/LDiOGgp/O87wPGa0tDEH/bdaey6msY
kFlSZQXfK3ILAdprv51cMOAYNUo0uRHwlbrytVjqV9KAD4qg7P3vDy1V3ah2qkMcoGh3omxK6bTU
Dj+/qlPHISAgiDnutNnr3+cVVextTDqCEtyVPr8Lukr9o+9dmjQ9+6RSEaKJc/jRODt5h4j25FcK
qpykH4xY6UDIGxZ80usoa21K5Ip0OJ1cRViI1AxCBM0bo2WuHbvoczuy6ArqzHDe3aOdckbX69Qx
UlsvhxmkmiFcWGSVnRkda66TmaXnyza/n0pMFZI6/yKPX7Ygz8CTq7WUcACNfSXBKXu47VzZcXD/
bTRkawPwJXiJLDFwmslNgeMh4ZMdOSowzRyshgLvlPbauqUA/ETXTHqvxcBICHGjlnT1SLBdR4W7
ptu7bCHQFkBX3rGygcn8Ja61U/CdJdi7grKtYVCY571w3N/KI1LQyqO21Q0/nEFtlvIEuxazbV0n
QWmIaMw9LuQH3DVwHNa5hUjqgRbsFKtxktZ1rEzANxdMKLfsq4r0q63qOJj2h5Os7I4qJ5xSTuIh
8MyFerenb717NO93L9HH7z+BxwbHTHYYu2flFUr3HH90lIkEGekSQsbVXnZbL8pOG3eLAgGOdAeN
/EGA+GPKIk9N8qbeOIik557nh/H5O9J16pAgwUMZGfpUwmMMuDEciMku7ptmZGK+VoR6+BJWOgb1
gNJ54R8rp+4cI/9jfxmqevUCbf3iBQofr3bie5YBknABWnM0qkNFSfCxY933A4kKBmYR+iReCrAx
67z5OUYkCvIPh3fReFAsse95RrxAQzTQb/FhHF4du57stBdre1B68pRiBYvmxqniWtDs6CwUhB3n
8hheDC5XWm6/BlUAD7VRUIMqZ3LVejyt1jgHnyw2Z1QrcdqPzhOQbsqrGCbQw2svDBQgheDla+eP
rMhBpf//LBEyffBisItdyEtDXDH+7v5L5YKzN5NuwIRRat6JBkvCJ/sfI6pV3mIqP7fqKWASba7K
R5ETtk0DBiv53N9k3N3dYGcyEOuuuMyaSpXRGMd8PIvZxq34gmOqOBBznHKq0Gtb0aAruqi5fbgN
jTvOA2R6waZ2uv9mOxxxuJwJfQV03YawKlv7Ah91iamc3wbOJFlAY4fjEgGO44cjW5hAiuVa47vS
734nOMM7uZLY5VXSw5NdpYpR8U4iUIGgal3NoTVXlgtoyCeGv78rFpE2+e76XCj0gvg26z8OaD/i
8BoIt9JAJbPQUgoCF3rgW5w+k/YvgluNmvpzNp521xrzVzQccbe3VaSPbmEpHnI202vGT7xu5gyT
TANnghMSphPwIRZJFI3owLYF+ULhRsrm3ga4wCeRAVCxJqhZaibssfW4m8BDWxQNbuk5mWddbGhf
avrkI7byGma/ZSv045K3oW6J9PsorjMtDSIqOzdbWI0NYw97soHyjuC0/riBqW78nAWABSJNoSBs
2Z9/0u8rqen6+3bO2R05D8FaSuvRPALAurGQ0gwFwVLv5ClYtpps6tVT/oFoDXZIIjKccbOS208Q
MzsKRCdMpSZiQjlB2qAXfbH8vTSRUkdkM+1CpxUzLX0EF45y8DFP53INlV2LFQmBCTVyrKQYzn9W
YxAixmDUny84/mii0lrV6yI/bmqyl4VJ+1u3ADFvNj65fZa5d/YrMcabTBYuCuz4aVIfEh0lIUEO
VgzvnUduBT5fA0QzB6/YFXNXZ9aGVblBmvm0IWwIfsnxXxO/mhPWptHrQnvJpY3Fwrl0Z2rVL3U8
QEzsrCNT8Vs0ix4E2R+w8RBOxbub5+hxb7MmRVhnSTg5NZZwnDMDe1YotKaI4oP19LGt97rDY1PX
zOaB5xlcpk/XhtvWbwiAhUtgQPo2vizt0acmffUndcyGRDmPhE+Ir0wXLiDKAmgulh7Hd6lNxgaj
PlG8MRAFOHbIqAP3blafrIXfsr67kZeNxtoyr7wBfOcmrBsQ/S15z7Qe5mVuktD674whayqfh8Pw
FPfvTyVdGFwmssKCE0A1MaXrEUDUfRZrjFffI4WnW9gx1wB3QqEDz0tBdIAi2uDljKNqLS/SFtl+
fVWPXz9o5MpSmgQuS2ZujotRRzPwiumz2zZ+auY7rq2gAFMSVyFcn7lsg9XonccCvdRlBwPHhkrR
EfB63ZD8AdN9Jo+/JDct2DexjMm1TWYfpbJlEOxGAmiJ70iuannQQ91R+7jqzQ2saBuAevWljqkX
czIVNEPBK6MgSVLORSF61P/Mide8Ud5cg1/BrMH2shOiIfBF2OqCVFN6gLzbV644aYDvNbN6c05F
6bnBXn8tGHZINgZTMueASsm7rLH61k0aYy09YC8y/VdSW2dQZ+nhjqNox7nxBMR7QjTpjGHfrjrh
qsVKrS/5q3udQUN73H4tL8UZGMbRdwQL7PzY5yyxJEi0bNNx8KxfxbPJ5HP2twUjVOqzXJJ3dEtk
4XgA7XyiSKff948LAUfp+Rw0VTNVtZGLm8ojUBR/YnxBfLk7xYOPl/J2+tiziprTmTsqIXWXxuzk
RQ2CU3EgxqH4M4T55izZt1k1L/nrrWmcEEFARskksk61HRJo9GJi4bx+2wcHn+FkR22aC8a7hkiC
ltut82z34lkxZCl/htKd7zcafFXySf++6aPA4VgxkzxQ4RcQsJjGUl/4QsfSWLE+RKvlKej8ddOg
//rbzlEUkkpsJblnYIigGknaT5vfvAOtJ8uKD9PL7Db6Ca8JFh2Q4KmQpqA7dd7lv3O9xtoYWBAh
XUjUtAAPYqkO8PXIocn4v8ISRUecnKy8JMhrxhekkLpA2D/wWR2eSxz+G42a00AZYWdpYyKEdnXd
E/w72GWfNM4ZU4qpOvhzszcg0lGgmiDbJivx6HVKoOV12VGXMwj35vlfRr7byuGHenyi+PBwvdpP
LjFD5GLcWAqMemqZgFmKtlPQTmS/fG8XOsH4j2JlSoaQCK5C9tSaAXD/ZzQuCGRDh3EZcBl8PIes
Jz29+Ssju7QhQ+c2d5jptAsbXh444162ltmEbJJP0ndlN6lJRIWiRbr74Uqv77/Ppuu3WUEfZ/lA
0tAVhHZ4xFAczl5SqeHxwtSf1recdDT/4jrC1yTLsKz/RqXWe96heNcHGUoJnT9e3sOUcFS5Qhpv
4OOdrHnmWVTk7t+e2saOn4/P6NTtpZC6wpGutyN/f/kduu3gL4tT7yLWU98NjmkTtUPeVSlvudJu
Q+Aw2iAvxU1FK99t2saHoDT51/oHTv7UiuS4uAMjNMNzT8VEESFDtQaBSbGvEwza4ls3vOGOoCkO
UdI8kJxwvs3mQRogLGZEKKejuwnSJyLk1UfoNZ0dsRwGDT6YqYDBhfoy2Ka4azOIwMFFG5xFZZ1B
NkSZohJz/kTcabQc1L5WV3gokScK1L/NeyoQrVJmvWEOCusoZgv6wP0Ju3ukDLSM00y4QSLuLD8b
rq2iEZVy1FL23ahO/o3HJsnhbdlFe+o+tB118q0Xbi6FyKpICL2dqGjJq4eKgLjQ7PjEuGGsJ4NL
dBstjEsABsDfKaMXS9qvreBAJSZVBxMFQiUy9n6rL8q8t6Io12uMWl7t2+sLcOppwG5w1lmdNUjo
aq/jHSp1zKaQ800/I2N5MOHkr4nqGOsPxBgm038pxSpxzcxiyf1KBLd9Eild5x5YGNeMAQ0gCCfI
DCgC7BSCF+Qu2HfGew5GZaU5YmZ1utL/Q0+Iu0XNaSjugdtjHBwmSQVM+5JArmquEw0DL0DZ/c4q
RqmwEyTRbjdP95B0qxc6AHJdoVMCS6m6jOzbGoDwSnLghRAB47qDvY6r1VtyClmtY1JpKslLfcS3
kwH6evPjEDjInYArgcdrkFiP6ip/3TQyiIMDPq/EgNEM7lnT75BZKtCXK62tZB2zF3wRHu/hdtvd
uotWbnv7dlq7cjp3AXeVWuHTDz8TI5FAuTkhgvEG8f9xL4D+jLFYBFsi3wClKUc4F8fzeSAAPUW+
JZx2VuCLuMon4V3GQo7u4hIdf1aj7oUPWtEGDW44do+w85trWzDGb4rz4SZbUdAhsvkTIOwHcgND
/AbRX/Y0LjVzFo2GjsXcZWnE9pPAQgAwXJgEVtVHJXOsUyFusT+OlSL+lpMHW7h9DbAT7slj9Njj
Ykw0swA1icZIUb38SMs9vRHk6X1TRYbmN/eglS92UGVUEfzmG756iXC0BUYqQQkpO1rqhFgED81J
Vb3SRA1JW3j+wb/PvIhW5m9TlUhoEk80gDC9gK1Rn/tjtC8onAJUm8sTB37odKM1Kr4QS+G/FFvl
0jx4DgmQKGmQiask7JR3tPsPz4sTFLNwaRPl0mEsYJ29ojBBme+tCx/95FBUIcvPagzfgmxvb3D4
VlrPiFOlpZy5/HTuctrp3N5kyM3m+PT7pg07r/nU7K+FEaqW7codsE62bpZGOXTxwT00AL1QlbV5
Yu3Sso1tl9H+fvSl6iZrA9bbBVdcWla24qpzr1qlS8AU6KwWDvSFRiPSpeXOCvKkEG5YDJ30TLJ2
Lrsxy1VCgrwazI6HQtTpdSWs4fDlcemE0LuAvT2meQP0xvzyPxhdUuiPtKxstAbUU7dSxoOpBgPo
uXkhDL8bKt0UmtDAxD7sPJatQlFo8sZ13pCoBnoB3PxS0ZjUJfmDMekvbb5AnoVKJx+gwfA/ml1W
+PDcxUZw4hyZc59B4YfydNkrMcY0RHW1yel9WMDfTUOJJf+XWVRiKd2cqw+8S/K5sJaYq8UfTqM3
HjbqiySufk7XdV6lgEXNkqZDUf6yMIB7r3L1QX6Bj/M3Vhx1w3yqgIsOuESLpiKjhPVZxEfx3Bmz
5SfjhEWEGAnren9pp67cTrWScjs1uy7fbNU/2H3aTithKKOhB3Alle10AMir7ehLnu/qSEWMCLPC
3pJsM2dt83wgJo5zadktr1wC0t1Y/rAatwZlKsexwvwK0y6/bSotxAUOMcwXYZk9hPFFLtZpkGlr
aTxBlUA3PxEHrK9myehWTkjbTxgbQwvY4V/KEILhAHbg57eL+fUnV48sEKkCB1lnh0lovF1Qxa7X
iBOds0MBCAQmFToFpiYuj2yIICSivTYstzZ2Vxgj7ety8SoQ+YeYDdcwkFy1/snQ/7D74eemshns
dgIevU6XyDREa0pxKiiQgwJ0Vi2TLWowGCvfk28eN3N7evy4ZqBqRQZwtOGSV8wprWK1rZr/QsN7
dCw4tXeQ6gsorbaItvVBOvcGM1dVFFOxrvi6TYT+msEHyQrVA5F/amnawr4blEogYctt6cClVs6N
62+UFh///AH8n0YTifnLaB6xiGDJPW7fsfLOZv7IjyMYDzoQgxLOSqP06qNmj2OVfbSHxQsumHOi
GYR8HltBZSoWMy7ryvDH1bxnjGhlfqAmK2qGGAZOPVAIiCR2/usM86KlD2xR3dQABkb7qJit7GQx
m6nh0qq+0QTXxorrskj1BrAazW9ZS01IK4pYUHzGJbUU7QTtLMY+/XEgSZYfHpBkkGZ6loqjZUo5
pSKaLW19KTt3+kN0qlutLzSFuqmprOzq0dSB2lffnT1l3e4ICyNfR4l+NTrO4luOSzqkwwJPy5NB
6+FvNoigvda+bjXSX5UrNj8PP/AbPLUAt7teoLKaaiAqR03lAQKpaFo1E0074G+1Ja3WakRcXXdQ
xuYP+R9PIF6HebpVhUa1mYQNSIYKtRP1AuM/MHFT8ALsoL1a1svV1Tz+LHhssb1F7dXQRvZU8e95
vARw78PeK8cc3bgaWF1ZNxAqdb9o/NryxVorBxIZUoL0//AqOW362MXTFHYDIT+Ybpw3GRosAezB
1KfxEQgOGY567ibE1shPVxeX/A8wgjgE6RnHrXZQQy9M68ZNNx1dXxMzxrRan9o1zBQCA2aXE/vX
CjQaL4nG032/xqU9xKYg7moDWuXXH9oxFO2Vev1jdjEpT7XK+UuZ/uoEzLD44Nvtt3oRodNgO3Gy
cIDwUs7CrKrVI36eLw21nqNX1ecnGm7Lmr/tPJmbAs8s3XpD6/QyrslNyuR6e9VD4qBinX/075+L
jrZ7esDjSvnLvtwCx3A8p2fhn4eoGfQKtj6A7Y/AUe774wLNkMdWxT2qBrIemaKvBJSYkglE4yx9
QrMR4NrKm2PtGdt3tZsBL+WjfnHEYr5DZUBOC8LOwaT467ApIw/FCKjvydLdjh/5NScWjnpJlsCw
0iuzgrC+RRqif6Z8kv7Gejqk1uCTpkY+VuNvJ2wzTGdLGpqjGght+cTzB0X81BxCv8yNe4NH3KQL
50Q4m2rdqOUet6USKgmK7gmwiW3FrlyxoyUTIsUnaMoVl1qZfRrN5SP+dXxvqa9uLsvj35E0l4r3
pZg2x0n/r421MG6A0KGQZtuqstD2+tlgClqCOKGMaLFIqhQjVg4ggI1gNlX8QNeTSCjkJ+uEDzPe
XTjEUFdNFtSc0SNDWjCTgOE16dPVG479//CLYSd8gqxNdpSpubcSjTiD/ZovMe9vbjC8fpITwuyF
3tXBlTob8jlT0VhdzEZR3ZtCkt2Q7AbAQ5qmtMuX4w7TeuOhzpQJmiU0gDKmlg1wgb7esJmXiY1Y
iCBMpfwTc9ww8g/LVZqxZWnJcWXD7HwuCSHEAJo+hcRhMFkv8aFu8dnmTRS0FbB4nR+y7mtjJ7bk
PQm1TQyhaRaqW4yRvlKG6S+dgnK7b/QgUpY+jWtcmnnB3gyUwFwrWUejrZQ22kh7NuEsMswO+gCj
u17jjNQuIUgSv1Q6QfSHndM05ARwWEmXVnQ6cKZy4uoiUrkcuDTslNdgORixK92axdRiGqTuhJiC
qaeLL7rgXkL5wglGPeiNZwtOnQae9dwGcG0ikUq7Y2Ze1V1rjuIQS7HIvlI7FI91mUaM9QW0gc+j
QM6idj0ENoctaYAD9tLefCZyxrwAq/RB/86x62rvWOLUbNKMLo3KzbpPGQ2uMQHWwZEu5Fc2aDny
aItMLrlPE6+0YkPjEw1591baHdLWxCEdxRCf+ig0DbF+L+fjaFJNQcIhK5aVI0BtX7qbzSDG3PXU
F/8hQ/TXGSYtcvDTlQiuQI0wg1wAuxr0TFSz8bslolK8+qmkNpvIao1u6TgbuflcRhjcuTW3PQEs
SR434to3H7DvHN9/4+Zql/uXDmHWu4gJHo6HBG26Jk1FxR37Z7mANGV949fzs8EmTSdq2HpJHkat
Ohtw23p0sljKMLtiJklnLJWx2ZLdYtv0lSuTKv2VMzQlV6LqqFh7w6fzHBRgiKYHQblHl44dc1vf
vgBgX1NRi5vCoIhznNzr4MQjGVaEyxrlmPYbU3lVCGj8m431KyL1ZnVMv2QjMR7qpYqx6qHaUDqc
/wPQ4qcf9+ZKWh21fzFV681E03AkXwt0TKumNHahdlK3NxmNz0ESNp9cHUOqSLu4EZLLW/jZjtTU
bdEQdo2xpKqpMZqCW4uzR3aNpXSvpjN3nMnp7V+GcMLnCwn0mBn2K/X3nFlFvzIXhh+MC426lamm
0dJNJika9yHzz6RBlaKrEnHJfnXwr7D9CBTKU3SBPHQCMskgET19PiF/BcYH+s6EZar8OUiqg8Lz
PmalXs7KsPpGdqZuExIqSEekhzkul8TOX4Isp2jcBw9tsKEiUuH/VXCLW9q+XmX5Iky2C5lwTiLZ
wnwa5cpSsq+4j870IShiJFjIx3CMMOChdC0McuO1x4P68yrSSRrY+IsanPU050ieqKaSnBHSlPNm
wbYTNzJnt0PRrf134r7s81KRsk6clH/bjQv61s/gKyR7LPqUiRMQxWZH47otJcmiU4NmkBEpg8q0
XIgZcvY2qL4JWKM1PguNaKHhs2hiqDI5jfJJlmcA4KZTWcRWSv9CUGZ5/qwVKcwlVdRosfw8e61S
0uVzTldkkdslDSj86JOk5Jrzqjr49Md3swyKto1UdOGsFBMU6FJ/1TYcHaRd3lxtZrYk4HoMzWJU
4v3kOZlFbwwvrQbppJDK0QdzdCK4Qiuvb5rX0dPr6hNmmoIRtWZhv6Z1obzmidnAOxyNiIZ6d7RC
2b6wEHk8btNaUSxL0/Zc0dve9nlG9iQjtSFcXwoAjLUoz0GiM7JURQ+ADKzFy54TClSCGxilQns6
Nl/DqKYLNLnyWww4bIeowL3TteR9ZxbFcxzDaWnAgRPUKrYSFdFMMMAYpvZ0Kmaow/ZtNieuzIKF
MffFV+O9XMP8hbnyUrXdladz6l2IHM/yfY/Y9IH/z05wpOmfXlFXLkYQCBBNrO2v2GoX0/ynR/lq
JUyvVQSQLyjHE0RhmHvcnrRA3DaPllmR3DTt3dUE0WmLE+6qAbUobQjQZJ0gCfqpKR0FkdbgbkzQ
0szVtduWsuZMOXmlADYkJSwwmdSnxrbouNuXouZyKgxYgv9/V2c/+clKRiWQWSkBrfZAmH68VwoN
Jq15vkdJ8tb+k2T29R89DGd3Bgu8i+8Jp1zTOxHcQmODLckQKwoMdOZzRPqFf2KNHOCPsER/yNd1
CWhaI1+lwAUtHyYIiF7m+HwTqDEWWKrmWRsuP+l019tXcGG7+vYBjF1pPhmIpbekqvJyYtlABi3U
EyEkV+vF0JMeIYJ4Puu0POzUg74f5tbKQhTjG9h46p90PTU8KRdTsTApoOKQF99PuTmMJjF9hTx1
do8+mFth1R9fjTRf6Rc+dj7pAFpuBXPY5x9Kkzlza5095z7QoB9rF1/5KdiOGQLW68dTPVdfLvKd
oehpWsPYJXkR1F+gZgMywKdaMjRGDTYdOFGbio7z2jjRHG+gX3OL59GOIiVDS1QbcIMHETRVgaDS
+7wNSjwob7HteskSA8YRAgSXKPd95BPKJ8+b9Byx3OooWONwseYCrdS5PklFQvBUvf9P2qN448aZ
oONRxpmA1sj38N/4fNea9QbZIwRpF0NBII1SPWnW8xcAzQ4jed7o8TQrvYJ+jkioKs6zqzsiqFUR
J1bMPbvtQDRWZlO65fAl/sEw00wImXMIeBFIz12ZhzVxGqg26n84Nga3ndHPokTwb+p8De8sc/KK
GucNyLZyNCpX2g5IRqiCKMKpoaYDpAC8uC1wqHUEV6a1Lw+gfqW2Cx3Vrx9iwN4KsmxAoV8eGgpT
wjYf9ugEQXbVLX2kO+U1boeyUZqkwZRn/lJuUCSH3cWiESxTmPXDmeN5+EyPoUAsYUyj4PtCaoeh
JbcGD21ttbEqNB7NQwq6E7f24p/etN3Z4+Thk2BgyEVHhgRiMGvJfkJFPn0cz0h2b5QSUaf1mKd/
84HxbWTUF58FRXjjtVmIixe2aN3TZjojLFQ4BifmyN6c3sGBkWt9esCGrAjRoSXoEP3JNStGWW1M
3kvbxxSeVvzjzcCWUpMwYdE88/E6VKr9SM5MLcxGc+9V1+i7upMBeaiHYVseC3EjgZvtebiikEIp
QxHaeaJkHuuDG4IprqIQkcJmVuFsP7Y43fHNFTxI12DBUZ//sjzoujyWGGV/7uYEyxenBTowEGAO
Dpz9FqdhXfb750CpYNkmyPISOwSNtI36zjzuAyOmzggZNdql+k2mlA17MgR+JIIe+i4Q8auWtjKo
t130KfhTa28WIUhyQJ4BeQzzZ3cZZx985l+JVO/Os7XYXKs641pnScKoThZiojy1vRUEQMjPSiGJ
9pypuEAU10LmQ+LALZTs5kKkOo2aqnCBGCFvfSgEBAR5yVdzJwHnSq3yLrt3//YtWaPzMq7nJMZP
Xt/ePhsee14Aw7GFHbcxRaAgQLcO6RxHQMhgjPQM0V0ZSQ9xKFVscxgBLz82CnzF0K91v559EjB9
JDnYalXXI4Rz5TUtWKTqWK7l2sxzDGME8OKTsKk82y2LiYuA3pay5nlGq01F+NWQ1zw1Fl9UlGCW
nWCXx2YXfw22+Nd6efbuIxwHlQzUF50quloMLUwWOpz61uIfGUCXN+59tQf3GNtESkOPinrz+imy
gAvxaGwEvxD+Vz93f/jMbBa2e6jY2nsQtZlZETYIFerWk3VSYpo0l9aqZZsV8smbPxKpwI/aV1Xu
7fMKkuNLJ5RsrAUUDXAv1I8F4GtIt2XP//sVobKoiN9edjDQOB5vzK1BSqCq46y4N4b7prbG6aG/
fZ5U1xH5fFchF7BZX/n56rzPjTftoVShasROWchNCfzChRvNXfFR9LPYge8ZzVloUk5RIxMgDUf2
5Haf2HH6llXcgfdEs4BFhhVvsBZJNzbQdY/rG06JFh+TJkYNzrO5oH6W9wC0hRjTlUxJ9785BdVn
cwLgu4OeVDaQhI/sg7XrNkVUL7gc/TiIinTdf0gfQIyhQW6RnSotoF2WSIbmLTxehVIRtBWaUjvd
h7I+6SdNBq9nkxlyXgtuttLwGIfgAddq7GiL4/FZMTniQkpYCBXcdeNKIH35PAAYXaGO46bpwWou
9TaaeYcHBYJDMu62S/RFvF5ZCu5yznL2b/v14UN29mu6QxoeV0QcjEwAvktxbTI7PxU7QAJfyiWP
eDnD3E6du8eCD+dtzcnLQcSxYHRcjsLAgrXsUbbLu9jUXeDBuX2RSiUiWAOUm8NmGXWxJvuOvhMi
xN3ZsvAMjbGfbGail5+7tSFBwq/z4QBf8cTVVmPwEZUmxzCFsrvwP6kJN9xvV2r4M9TjRI0yGDeg
mpyHS0knmWttdnOKK86Bg2WL8HDV+7pba01AvYUjzeuyiVKUi6IW6s+Yl5gtKkPdoxki/fv7/Ifx
YAsl9i989xm6f1DrGX7r+j0ybRD8UCyc0d7/eehGjYmkw88esWSCl+S4X0NCynPi40RFcgm8pvNO
Ki8g349xYUA+PVAGDPTOm1mGLU/gyHeJSfAtJwKI6f17E8JOAQ/PT/vIrgQNdJrbPILLzB2JdIXh
8SVShrNEA2LZBkTJD1IcrKUfOv8OvvKn9HBzQfxnOHPawYS19UXQiNXLgjmFOvTdI0XS0EPUYhN0
aeuGToJkj3a8ODyQNxIhBZkrIaw60BqlS4YV7dJ030g9oXQ55x9TDfcPciCO8FyJkOTcouNtNjA+
b3oKotchcFQLcK4vmd+eCHQTLtdV8Uix8fT0iAU2L3kl0EiKnSoUVon994GqXLIqn8MXFlrop1JY
mILodT9PyEIyTVIuevN4aDzv35oCEfeGS5sONwsWUUCwu8pQMxMfb/SxJmhw2C01q3KTIxm8tIKa
+ETmcmQASLtnZN7lNUVPq3vOWyNF5Ljy2ARNII/iOG8KBRrwnCIWglltkiWSHO3O3f6U7C4Iv56O
gpnsEdZkHpGUYlqFb4EEDmXrUubAsjz5nOvFblUUxsnYeuMDEw1ovtW80nZ4muAzeylfAt8Vvi78
ZNqqwsyHsrI7scuKZXp7ChA77coJ20SiBCA1TwUtMG6bpFP6ZYBDXww03mpoYHGo3cSpPRnV6QiW
J1AjWUX4X9t7NdE4334vacvNbma5H1khBgDAapR7X0XlycCN/nOgoXaPMy7CIBjx5UAX4ZUZdRwP
7ODV/iCyowHp9uF/jhQjNUtzu4mIr7Luqcem5HXI96PHjqz6xYhfIT5Pd8zTsopHSoDNibll/pjb
GqKtDZFv0OFRPxcNIqlKZMxIBeGT4zlMOUp/ShIrGoorsLM5HLcxw/hRmMeOvymr8qCUX/jFj8+7
IALh6lwpNtGOSotZXz4J/BWqqBx3S0oDBNWUKBS5tFb/2PbBQJYMJi1yxhR84WEqmiRJmsq2ltCg
VsiREg4d/3kP2s1846kvGllbfnHkmVsWrtw2gNDezWAr81hcxhTkKDhejtZhRPE0LVzCL8GC5gi0
rE6xYu7IJ0xVVY7pVUeEIC19kjhatUv/mt+8oj7Y5TjrOei5rprK9p/Nlez+Fd9eGbcCVhZxDfk9
5LjVwenbGUh70T5eCJtFkidC6b51Bj6q6Ptj0MLCrY7DAwWezBBJQzoDpNUBrd7u7ZRKjOGCbCOv
96VSgvxVPdxjlF1iWihWWwpfmRmdQu2ZHmo9EYi9VjBuoTEZ1oyDfhtA7h88O4sQuRA1BWTtDN4w
mspiTbPtLFfOmOsy+vjsvQ6jNT/kfwS4i1lL22l24eTzq/TLMM8anccsb95J61qD5SLASI9M70Mj
bLDiFaQ9Y+YybZUOHO/FJ7S9LydbaQFJqYC+Wr4XggMc6CLp/nJxh/lJC5rAHXXsktJoHYkuguRx
480pgDZJciJldmMogBswbsm5aD/L195/k7dSpQ5krXvnKpDxZLX2B68xl05jCGymTx+PRNhFnIun
EEAQwSPtt/044nwInrnDEPXokIl7OXko9j7vEybzZ5yAsChhIVJUJOdcvSlAyuU9DcwPknVu7vzO
J8ZCj2tfdHhVyS9G4ocWOPBbeFbryXQ13SZV402Z4HbvOSMIzLIB54UppxM6+ETsNLRjuWkqSoCT
VBdRmZ60OgJBpfWmnccd5We5VbrjPgLFz5G+t+eroouGqY5b6oBasTjoN9cfagBDwEllPl49BYbt
1qYsfzoAG3BOwqyWqeZR+vhwLRw7Jycbp/zkaiDJFIpI18srLXwahIEPqn0Kt8HCfLWNgg1hr1DX
46CrNqmKWRjESSH2aPuEz55bEWnm8QhlolJ+SdNyeA5RDcOo+jlbXrFgKZJ1fOQaeuO1s8xuiN8X
QM2gSycSbh+SyMVoJdPBh/brIfAWvLCLGcA49Mb+U+mSPc9192+FPakJy4nuWkTI5qgelmyiFgBm
2JbStwgann/nSfMeWC7KMt4abXgFKUmH83rzTS4ZSB+xZLCYu4kS1L98BfS+ec/aVRjsEVl/xoCb
H3w6YWq8FSs9aabDU+ccZnZKDPfBjfgnMsV3F6svR9AiEOMicTJ+rgG2MKksbWBzz4km8UmmOhae
oRf2r1jeu9IPz4djTG0wez+70KUg4vMgRdaCX0njYP4L3GwsYJwwFYSluzYAl8ORs7gr/SkR+YgV
H3IkXGzwaT6RzOqZIiulS7DR2Inl7Za+8NIKWwx2M6c7u/kBsELl+Yam4aKKnHZW3a35WdyKlR2M
HwHJb6EKcwUldcvKZccrMSyl/ZUu+tFIbU+wG4GQ7AMFQh4WRAhPwLzayKbmzt9zW79F2SqbyrE1
GaO70uvaD65D6m6Ptx1tnM7M+B8PJl40fd06Hk8bJk9F0unuO11mItnY98iRQN/d2hCpd68Grjlb
YAvfE53z2Bg1BkxrgrbMfVAFsMhpQ36VDqy4KxVXO6sOlkIYzSCMxlbkNMKVeLK1TI7C4GV3TnAa
Wa6I5bbgI/IJl66KxgJJ2uH4cTkcf96WKWctn5y4wIHFOI20tIp/KbCGjKn+dHoPWMV3uObuaQXE
GLqXJQUC0Y8CIVRW1PSV9jhxgpM37fkv/g37sfxYOb3VsZROJ72AMx9zrXl3Sbtxk0zNVaRQc5mn
DwM2sAZi5F0a5N026XJXLuGeuEsKEL6xq9i42xJKC0lVRTmGwa6bbI7H5jRKxvNix9ez8rpKTldf
9cGV/rmMCQVEWCq4CNQUKvXmZ84PcZImFYsmZPrtT0vMEwpYMLoflLV1zUPHTrddr0tlzO3lU0Aw
4pFNQjcQAJRhn4FbUptoCH25+8S9em4jkxRsRnUPwnyXgWVQ2qozGQZsZ5Ni08w4oyNLn/7vFjw7
h4+yCYT/5mhZyNdzgGRXqYZ7LiiXOwh73H+P/nVw8vRmRYoqCHmMkzfyinvmj7AMwcTTNw67NWL2
pqHxxE2z8sXGhgZaF+rP01nKt+urISmfZkPWF8odgh+cJGSwIaweZWbCp3vgFDqArUePH/nAeEZe
4VrcYuJ724VKxMeFxS+Zd9h1HVWW1cIYMH21m2Eo5AkeQ9Kl055o9cmjherX0mb3SijZaiV02YCo
OdxdP60R4iYPwUHXLK1XdRrpTLYpAZ/btHqPG8SdRyvQByKg68FQtO/wvV9GoHNLNjxIZW537TMF
pLbAr0tJzpzXfActbp4y0cf/E+MLu3PsMIz+MXhbmLZb0CmL1B/gSFErqqOkXQph3jIadFIvH3xs
MgvreJ1TAzXyzhUeppGQUq2vuhnlcS7x+aEKY/dbIjBxZIL/ex/s2qqHcUJzWttRjy+7tIvJJ6cL
zJw8CEKi/9KsKDPsHfqfBo0BFc2P/Y6UFmPEWig/Vwu418E38SirhAJF3MwdsYBC+TrC5uJauihE
5RAyblBcfm7kL7yNXdAUjodXbjqMurwHTp/cx/PM5tcCI2o57YEWG6SiAOIM3nB7rT7bO49UP6kH
xTFimhr8MLZByq1JQwGXD8JRf1+NMYhG1gDoHLrIsMsivA2/8IUpqRdYXHimb010fVJ6DE8MI4Jk
rpVuBUl06HEyJVOWSDLubyCDcbUKEzlV69inLII2fJCt+yKfNA8moseopuBIMtSEFOwnbQTVfPvx
vrHnXFCfhScIBGypBKD8GXNQgaJGrqWAIO9uRu/HQrGVkH+qM4J5HxI4Ue9IwIpHtlsyrPkcVE+h
viVlzVQ3vtaKEP5RSXCnr+vpKbB5K3cJPBm/um9ZWYGeSA1e9qV5Gw+1op6MQlcS0RziJZJwK1MU
vQ3ieV4fqpbLX8DvqFFg/0wa/8tbHcy46fU7XmJ5v5MVcMrdrcvI3SGS7qO93LODVhjoeXNOKBKN
DnOA6x6Om0IN3GT0bIuPTQRAXLOywwVy5/VSeMAfos6nP2pqrAhz3olK3l6O9OV0LRTYcHwCgjmp
bIEZwOls970EEprFvgakiqOki2gfpqOv72Widwt7HU6f+KbECLUoAD9YayJO/Bbdr7DheF+2iQLA
xQr2pITx0Nz3jVefghHJ94aKzmPs+8PpIgcttVx7cqUgfewhPlBGjW18hLbhgWRvyBrEFtAzfnty
C2CyiRQI19axQvPJ1Ql6RVW8ITBn+4uUhQf9ZsDB/M6rp6RxoNd3j8lSA4EkhIbNbBxs3OCYq28f
MxcZ7OqB9z+/8/mZuZ0f4EHH8x/WD6P0cTKcxI2d7B0UOg2yU1p5QtAp11poAlnBKY1XCvWPerzo
7XWcfutGgBJpqUp/mnHaTt1R1CcN6pzk2zjrUcMgOdF9yHc2FLDRMEuAZJG8L9NgIMiOom6He67r
oK7tGfUW0x1+hX3xSexHuicoxstNiDVfDjHC1T2GLptFw82VakMMz/mpk4K6KlXQeAtnZRVtoCk2
GAig7ZJrPn5X0sQmU+NS9XBLavFJuZM8HaQPB/rDlgnwH69DD0ekrn7bFMDfeDJPd+4v5oxeS5HJ
bu8b9LXK1B7hBGYcdDPh0mgdOPExSB9LBIP9moNuF+lJYlejixo7h6fpQlYXcLsMWTv06DPMxMRZ
4MM5HWTQVujY9/NWVrJq/ObKwOxZYo+8InO0MHkc1vxTuvVBvea5qIIcTD0zdM85yWP7ZRLMEubY
iZoFYbnpkLa4TCVOSeOIhCjTBcWo9UHVFlQ0ODoGpBzX29zeME1c5tfoTkazhHDZ3MnyfSCTGP/d
2/YKn1q37w0d2iempdhisn3aQNpWgcv4IfuWF1wHZJ/jH4zMAmrG2UkTTZDxPTQGd4rMteBVBcMN
b9/CZ8+WgHnlgBq3w9FHG6qW4w2YlTMPfr2ox3J6q2isGNghLpJGBhuDZRgaL89FLrVQTS0OwvFi
SRhvolpIEFYfELyHL0M46UDuNUGkEmOjrk5Ca+OuCRfO9myRzlYTy1Ndpvoo8ZkfSzjUGINoFtBt
BNWfBtlTQUcAQnFosSsRGVv1QfWrK13A+j3fvFBE6b/2Mga8brDbMpNtftiBS1NjdPP42I+ZrlNc
KPmWfyEU7LigRR5OsDimP0/83jeayvT2Vx08vjhZ14cwUOHrfhEXdjiK52Sl0HXbChavU3GKCVsX
BC21367+B3N2KUQVLQcXHa7ucIZXSG1g+Kp/7kornBsYQWWQ2pafy42yVtG1pCTtFHajstGcyjPv
OCC6JP1wIP1Tn4CrOSf94SZnD3nV1ibmmgeFUBE5pDIDgqGrzBVyVjG8hv1A8Vdf94v0dMV2HcRH
ML8wSxyGq/TIwWnbkNC6fAVvxmJU0yP9wfk/9d/QCHE1MpPYIolCFCVTZEgy1usMxNFiQac/qrIz
qPoBw5sKSxkD288r4uoCkSSMyeh4TAoDKmHTeq7atNqhpgRFZvwWtPK/K9npfWl45UHBc/L941QS
+Z6Xuh8+pMWv7L4t8CfkYLwIhUulg5dAYSEn7NXLLQjQuO45+xzwyEsrCFCSYtJWSJ77CpXZ2/B9
IuPBzTXbwV2OJ4Un4geLKvso+iKULQKxt69pmTr5HCqomxxHzgrHnQ4n5mxMvzjG8If7x9z+JxT3
yhlx0pjYKGyByN8ej6MWkmZdVc5OexyEAGy0itACGLin+eorV/o3MKT/Y5BCnRqkzSFmjWN+hsnJ
+F5EXCDZlBt7Je0nrr/fMOgSDJVW9+U0makEzMH+7KUVpmBxtssF7zQoc6YCK1H+IWzDn6NOQxxs
I8Inucm/nqyru+RmDKplDOnZBf396tXisgq45PNtt7OjGWKRHC+TTnOlsKLj3soGcBZTpZY1M5jd
o3IXptRZ+gfFWG140zMK4D3iMjWNUrQnkQu7TpNGygqVKRVlbBjeWmKYUhHqYXTQSGLXS6MX45dh
AQAPscU2xSHShfbMQb8XJnqCO9gNYZ28OiNTyjf/LUpL8/d11jcIlwLiwyDOVaqcIGu2l2dPO4xq
AYqIdeavVhfAIxfNtIxKA8ZRwPKbpmc7Z9LJrg8W9+eJm2eAwrBmCPCMiazFPYV6oZBMet2saBLo
baLPVNRTQl3Q5EGbOJbh/UdWp6j1qSdMGaw81hlUBYjijbL8yIerLZVq87DlhKg2Yi7WBY1u/ery
/OtuRHTB8YoThc5M0b/X4KZRCqgvfgoij/O7kBLIntlkpOwobb8XmCT8bnvEsVRNjTKEmD31uTbb
kFjq0RaKTBohhiJy77MXlnU5Fu2g23o/gig4pZSs44P2dTxkljA+bE5jIus7Ksk7K9BPUK4dev8m
EEymvBlnRY8iQKjQ64JxshL72NqW2AUGmyTrs+p0QN4vrEDibWyYkNKU/oVog9mvNq2ZLJvTJ5Cj
IXt+ewJrHHj8H68sumkxyINRpvctWtojM/iEEyP6oCX2a3j6pZyL0GrSs5taDhZU6AwnNM8SQYuD
zNh1hc4Z55jZ6t33FWcyLXZHaGcyr8YvjT8XHsa7L12uxVQlPDXITUER1gAdYymnLytWZXei1beg
kGyyPExWgVDLzggTBgDjuba5PoTrdE7IHsELVLcKqW9xrHmYufzPGJmI33bCO8GUmSsAOr8sXRdP
c/aAoNj4zdYzMeRGQNPlggsTgYU3fVJbrJWbgoEN68mf1W6Wy2e8kuwVcpAMJrLOJeqth0B6x/H7
l7RarFcv2dZaUsbivcxyRi2MSp9gwsZy6WH1GDacbCBK/Owd9xiI7X6S46jg5WnOANhN91Lm4hCm
OP9KU+J4KkRR8DFz5SM87FsieGAHrqzixPHN0LaEu/neBUgLX8obMLndSrCI3LvtS4y63aIv4QO0
cickCQo5EjhfjZ6sl3uMnrIzQ+sH9PX77hRqLl4vL52HrRWA7wnYFXkdB6uU6wM7eSNop788W7zg
/q8wAmvdArWQIiD8NmSlMKJH0bcsoLnaF6Q2/LH7WEwtIGmRbweN26nnp5BUkEcS4JR+xz6fvjDt
iIlGB5ZM/tbmt8a/jUHgS8xaXnbdhW6OdNQ3RQ6Wjau9wkDTbjXphhR1sSnujGXBlzR8l/vUkMc1
pWuKsqnBYg/G65xNQfovtCIeIWbpmmIT3eo7rkdvlq/qS+QV3ZTdeSxACILGJcGFKuJkZXmKDXpI
QeuWOGMFc1hD1sJoxMENbxp0NhEl52OAY+6yLd80mTTfjH9nK/Hmw+ukBNezobQ1nCTFPTtxyuw9
L/zQDwjVlOd2PxnZm5kHkzkc6UMLttWHnLDwC4njP6/3ClBud9Mxw267sOFrWxedEVgVQx0nC7Lv
bbBzQ37Xf11SznEn09oiqJDdBKIeh91EfY0F3omKaMaUsMVtmo0q0WJnWWNeRSBP5E6xX8LkiyAN
kEmsVPzJaAQcm1VF1ZosuBTpaZotjViwSfhwC4QZwnzGF0Rhr4wB3V9kY1/9bkSZTPsbVfq84E5d
LImc6gF2LmxDFSK8nnbff/vuUhk4ymjq5dlwVgia7rV7oq5N/fnAX/pc4/N6OOARE2ayAg79m8zF
g5QkCKsTZwlq0MGAYCz3KorMjIlRCfL9W6FFCOVl5kUKTm1bIqqztUorN6d83N15NR9m0CIjazxD
5Xy5LnQXXvjFY2NnJwUo5Bup5ZYhfGLQ5gArhZRv01ZV9PxfOGOpLirIp4RCwa0SKHhC25VuzZYQ
UJisXzM/hg3Kh6K2m2oBNRNvGFs9STFazp1IISNuTlLiW7SMUR03epwwwGeZ9l/N+8ms8rTSXJ2U
MF/T4+lX1hARkxJgV2+KfRbDOI2+rqLx+wOZzJTa9votLTtzpQJEQXRbzLGamIYqZluiKHHcqaGY
q/xkZumCQzB4XiLLn16xzBW2EV9Ieo2gZdpx6Qr4Pv+m/lm3sjtg7/4wxRS/N5RgvANoVYyeI3Jk
X6h5f70fdocw79FsFv8d3aaNmBzOtNkjoiRjj2/c73afn3nh6PtHXfDgutPisKunT+X5xqxkf79B
WEK1kat560kbrlMRq/PT93eCsXMexOn75RnbJ+yqsunTXpcnG4YQnrk04Syeyg4nwUidJ8GVMDaC
TDd2MCRwGD/LLY2zwroPyu41eR+hdBHCsvAMoIJnrYEnQKqnA0loeyYZPbE9i9+XRL37Jsv80GKt
ADB32PlSb8YAy9fxDACla0siZkFT+vXNgp1dJ3HylqaYhRJ+8aRS21st5cf8EXWgHI+hypHdTDjs
suAtpuDobyNNleNow5tOL9fjxdd9X98rerp+uSUOmKkVGHT/0+SgTl72iDVRU9s7X38m2oqxwNLg
UEZWLsn3LFWv1zA+11vDIBf8EpmtUdqIaZ9z6Z/hZS5SEqsux0FM1I1XLH+97sdyimjl0bgKeZ31
m2UXpi/kYiXaV0eXoRvYSXtkq+dA0jzHQLGLZC7mZggQE1v9zW9a1je80VBB7nmdlseaMtbp5Dqu
uITsTykm1VeiVJ3Aq+KWvMX2lRYE7eQ9LKfjE0tLo3jZRXriRVdqlcxzfFdnKFxrLPOIdFX148VV
NCSf3Bi5rbX2pAhD4vNarIvQqc3+awYfr3HfNmmoAI7uB3U7XQ2ozto09vhhRRE3qM6hPrV/3fBs
6ueLsZtHho4louxKhu/vDnnrSFidBuGJEL4zurWDnGTyXNsvFV4aPKHLhcm6QDET4MllTSO65SZb
uEIxlDWRvnpPTDkPKTye3G5yeWx/22UbNnG3TaWuAcRfLCKTUUwtbM9deZUSXP39H7QYAh3nLlIu
B/wFjA6Ejd6DJpkUmS599NK0a086eRZHyYpxp0floa8U1ta+u4fEYp4e+pZCwSz7Ihk5AhExkz6+
jIs1s6Arl/QurIx5lu7pMT5nA1RSAlwXn1qeQ/91EYVk0CIWOcQdcobm8xgd5j8ClhYdv/RBDOin
BvlQkYuromaWOXQfGKrtekT2xm9bxksspJ6Gp5b6KFM7Dpp81KPvx6u03+JcxdPNgtocw7vhXxkt
3dWo6v9egyfyb9ft3HtuDTsbzOsWPlMhrEjS6s43hDFENodSh6YNwqx2u7sUXwf0me6U8X4bfNQP
nWO7Pwd6pYfI3CR++/B+CauWlOldXkjvtvetS/oSHY9Jfjxhz/JoL6srQcY73SB/Ur2bl2QhCkkw
R7vkHFzt1pkKY8s0N+YhafjW4Ymi0if4mtaXQWLA8P4vVLhaIgsDctu/WdpDC4LYvrfEZVQJBGW8
B9/8s4qe0Ii2RtlvkfcKWOkbFyJ7/gKCwwTfMons1Ro0r0ucYLdIrwDxJffNpsurm44Bng80zM9A
HH8jolMLER3dp63CwhVYaf9RmZEVcy9WRgYwn2ahkRj/w4pDMmM20QDP1PSHHGzKfKXvscqByPm3
8ayb7CvXO/4PvdJTNkvkRSVRE8Eakhrr/VSasnIXyzO+KtEI7eZz40ZsYA7njt5JusAw4ooJTXAV
STqqsoOE554TRiMZiTOHrqt83prCAFllCkQgxDB+SKDiBef5NMjHtBJJz35qKyxYbEZ4Tnvkl3fz
qePAoDvwCrSUE9EZTTvIcIuzWy29yA9mZTCH0eKiJb9JgbKAAa4fjGCHxXEo26NqEChkVTffknyj
Qm2UdN0iJ0+KfxVXLV7AE8j9Hjz3sAx4bn74i566djGiR61CMddb4JTo/Wuq9mSQiee4/+7e1TnK
ukGB524/FT38N6JOPiWEyFWpYDjj1HXWrRnR4jIQt3JAJcAkRkbfSN8rnNCKba2mNsg6G/u8ARpj
YyqocVdd37Xx7Ae/mUq3ZNElgOE5cxJSI53eLBZhIIKr45n7VEjurPBkleKCb578RPpzd/Dnis/l
Ti4xPqXTNnFLg54o7f3NxVNQcyB2Wb79H9c4vHDCqv+e2oxBzf/BlLqbdrisQSikJdxJdH/WKa7O
I+nFDJGBe+DIqO9pFiRAaq4VA5o4pvvG0rNeiupCXiqhockscVYy7M40Oev4osxUa63q7iBrEPDj
hQsJrnQH5HXCALhA441skB9APZpeLld5pmITJU2ajboW3dqt/phGSSSyj+O02PcuE8ZZKYjpzcss
HxxgIJw12wcnb0z8re1Y6nL6wU+2I253hBoJf8XqAcyb+3UEqqpvLZK/n+xeO9h7FBgcOT+SUQkw
PAwtdFVFVBaiefGhxgFaXlYhH5ABPFyZtVBZmSNbpXfcfHCcQziCZPjDR+r8McESjsOmoOFFRXbJ
c0cVVShd8g/BUPBOagXhk0tLLaVkxNOvweoaY1kIROzczDPymtTs2nEhCT5vCBS8z87FEz9UmGIs
mzwAOIAECWw+lyBDYiiN6TUk29mUV1l/+Qy1m3myWbZsd1ZXwKUNXhelniLkKAwMLipdXPIRgjQ9
t79oSOEc0Nw5Niw2MhNFdCr6YoBUeu8KF4xPxvwElEtJOu8o+5pu/bOjOSgkZRQWbR5od1PBoLFe
BTfPvN5iXbQzAfoi8AVd2wEPT8TbsLhbLMmZW2JuWxYASLGR5//f6tPUvNRpChinn8nJtYtTC7XR
L8/iDrhO6HkGpvxCgWc7tSk3kHBlCYpiDGVSlCf8pGbxMXdyvaieQDm5VZQ6d+b3EaLUGa1vAjMA
osj0AqIcw6hnBRVL+07xOPJGzojHkv5WdARUqOrdlMiiE9ISrvNbLDmkX7kpXJ6FhjH1yKvnQmM1
Ov9+2cILIlIWWGh87BCs38TLRNLbtfgxnHH7j+vkyoW8iRUzOiNwqAb8EYaHY6vkP5GLqAkFKC3b
meaLMF6a0GD/wpDWaADbQdg5SAXKOdRyzTkQn3vXdAYto0Csizx9vZvdENQx3S+0ZxCdUsjFxlTG
Ts+w1Vj/xbB7t9jsm42mg29dn4Uh2cvarsuZ/krwPPTWXWpydo6rMRGFiUum+NBoAaFGI1w4r2md
zgXzEz4GfzOPMpLmFzfxhtj36xZn12ClaW4OK4ETpVwpbNWuo8/LGo45e9arN5igLRkfeQWnEzNt
sCAc2RfPkTq5wjnrhVD11US3JRUSu8ca/kzpna/JunRnDomsQ6A14AskqoH3psuVm8twDSWNBoz1
TAGjR9GBIaBWjif2OIrFkESzUeiqLuW0zq/BJr+y/qiZdyUFUUnmjhmItSjdZOQh4ZtEosCbxcRV
qGfDgIP5o0zeUedIHC2XesGhGcj2d5vovytsDRaRs5PY5p8eFOGc73Off+5tKswBuRCUJfVUGxMv
bbhjnj86TIU+BghG+OJvqs2nXAEAQJUVlz2+opqzDEDJsyS9m/ORsDDyIU7g3VYwmHMCHuwWKXbA
02st50xd3JkOkjLsTO5J0dEN3L3pa/sJ7p1h7FCI8zCiB8cJHAnA9mtFUq8MAwYakRM/TseQe0yB
iLiz7GyQuIsU3YXRgZN9MSvP9CRC5/boQu8ePuY2S0VJqi4UM2HIjRsYrAaX9rm8aFy8b/G6yejO
apGoQ5TBFvSL/3aB2XYqypnfQDF9aPXBNrJQjM8E1qZCT7saGkH4djBS8G8RylhbmAPJhpNMsJ7R
VAO+LQ49A6ISE7BvO7NxuMNPza7IcLbaFbWAwgGd8SAmsHxR9rbRQuhpboqbYKJoGiQAcABb9hvR
lCho7vNZ8lfkZUQGJ1udmUiOi4gbcZ5WWtagJPTRDZtiYc7jwPvwNKcamSCM5N1L96n1uWx2Ybz6
/KmR+EEvSrMH6aq4dzbHuXBTdIrdMXnG00PYkGr44lXg2czOtir57JEOLD3Oj01yboNoDUC26QCm
hh8UyWk8w+PkEHZI6aYDLdyvbG+6ARBwMjLPi8zNzHVQ4m2IiqsxaLkdJtDrOUbiIkYmj8quUA1+
EAp+tpBAa5CH63WSPVAJ0GRDtcJttDyRYPYvsW4jNznfGQGsYUAUQ1feQOD97B6MRB/tYBQ5Kui+
OoVFiE97+BgALzgHG4bjl6CIpQ1uJ0tz532mT7CIjAsSgc83fo/q23qnxqL6T20yksOoKLSztDDZ
Ey/3932egymzNSJA8B9yVApsQbOAz2RJS88MBEuODJtq5XqVcOI8uICjc1BgynHjPVYey2smCf9X
ExFxzpZPtEWLA2maBxTkQFgceKRPi9GSUfO03IkzlbwzCT8M8SWWOJlPnAuAHjQdg5zVM1bu18ql
sIOm6YSwNnQwpMVy5o9VBOMhouip9nVT8C+67o15rT8IsonMnSeH2pWE/FnldyxvSKmcP839sTNT
03wLvz/yQKFVM91p79Hd5yifU+KlYxsk2psw3QNBJiwbofoBDsyGcAeDEGNun/0SyM3KqGkKaGJK
CA/xzEUNmGYOEVD6M1z1GClNT54z0o1SIKSHM4C6Z5r31dC9Xe1XEBn5em3tPPkOfC68kSHklA0v
77kv8m9N0TG5JDFfwwhdsh9P9CoGwknLPk0u/JoH2BIQ5etO/ucWJaD3UtwGLW9chydlJD80KUvb
6jN4ZEKBqbJOzjwKBk+GAX/gS4fzkKqHXqq13l/e0Dy9oOngLBAyzIz28XvkCVopynIFmrBgGutB
Q/aG4JwZ6VIeroHf6ll2ihV0vWAX5O/SsDfLvatmE2ygb6NwXWw/Fszq+9cYpIi8jlVTrNhlM2b+
lJJEwdkUTASYnNfwh7B3wGUHLgX/60ub1tF2LEQIOCVqbwr6l1m85JVHp/EekOU22BWmayVkx0c6
vaHE3U3D2pc/5EWmftY1b8djKKjs3Im4hYkvspGXMVB9O+R3ylBDz/g+bSnZhn918yX+A7LpZxQb
EROHYtG2D9+3N1ZlmexgfDcpTHBB3OxgeQ3EPPfSzUXxCt5slGY3jf5FmKI2QtqIazAdgX5CShZU
uineZI74xOvXOZqVR/R/H23w9gJlmFHvD3df/hNwzuHYGYVtENhrbrQ6hhzLJlQ+pumqx/jIhEt9
/WBEBpb71t/xuD2StS80Hu1r12mOTzRaRLtUU7veS4KkMEOrkF6F36t/DvK7jhq9KxcSmq4mHrJ6
FylBU9eeONox1y5YoHbVflOWnBSImP6n/Sbnpw4dd+1hLXn1erLBnUgoS1OTFec3AWDOlnx2eg6X
UqksldI23AA+/IW9C/O5uKeAHRoFvAS5RDpN0/2jOVp17RWAASWdO+I/Od/W/WaBgZm/mXO3iJ6+
hWhgozzP9DbNvYIWdHF/7Z69PftTLQxxv92kHT81jaed/z5x2NBUrRcjLjdKEUGZUomj7H7vB9fI
IHc0Q3TarfbBSfq0/qjuv7OOsPHMqZtyytQ+VQzBdFOtJhqythwirmibFPVlIi1lXf8AU4Rt4+Ss
8GcD1Hn5A6OGOwQfXP1bijtW8yyaJaRRAj5EvRfpTAcu0PEa2JcNWgCeO212Dky4Qga9ZOVuPgLh
FwLDD8jv7uZxg+lkmv1SEqXkXKis6A929hs1hlHIqSn/cxIzdjHcBwWtr/p4+2wayxT7O+Hz3qSi
k5T4Jau1NMq9+3X+ADwHYBehncUCnYnSrcvimC6HN4SBTWJ+upECKxGNkLQ7UvHgSJlf9Gsw1J15
dEgwtNDK2/YwNvpyRnoigmESdA8G4Dezz/mgTG3+RIk4R/LpGAqhXU9DCz+zsftDQaeYONnHsphM
NQ4CZp7apA3psXy3EgIjLeZhjX8PUiDslRXTImf2yuuEw5ftrLq8u01l4kDqL/MXImrT6BOSQJBH
vI3WThSo1SPIamZT/pRBnZne3BeVOadO/v2VGOWtX1XjsJ2C/6EbUlcpFa5cz4VHIjXq6uCETnjD
0D7z1YW8rBZPsluLP/T6TiJM8Vbuf/hUKUyYvFqIoRWFzZqJjD3tnRTSvhWLLeTOvKRZt+A5zk5U
WiYvmRo9U0w26VubNLgVizR4leE0Yqc+r8Ryjwp9BsvpKQhwAfrSjuz/MnYX6I4yfYFCfovgVFrD
SFqjJM+WDMrGRQ+FyL5DEm22cz1pJs2tvqCKAh0IGatWYBjc0vhoov8Evlx9Aio+dYjD90Ntchap
/OWvUSfPuEYgdz6eQAM5VS/WnUYmvqSE51qGAglnL2I6egZAwL+/SxSvmR4IKZMKHSe78YIfslV5
QdK4JCYVWIfkCeYuEwPqG1IP54izcgJ8ma2Y28Qw5clfhajIg176eg42UC1RCXxgQbD1C6r12MJs
I+Enaa9WwQurcQjYhcKE4gVul3R/8sDO82Bnh0FRSt9CVpbG3axeICT+1Xm9YaOvoNKm9aeU4T98
brOuhfpBVsmaK25kcbPZr6MQZ2wTGNxKlhyBGAx40gBPOKQlHow0eaBf9Y3PUIxHCqCxg+fy6Nkf
BbD3llSAdtsKDr1AwY6jSxwXX9XNZTdYuVkcun/kFN6jvdR7aAtqw9gqkkvqPGwXd09scA95IZXZ
CKC/ufU+3o0kjytY+tmDw+E9FReijGdleG6Wy8yTm9/Y5exFFZb+nm+G2zpV5bLClBo8JsYwmQ0l
9HInQWbNjGOK5sn4/liVWXsqp8qNAcb0D3TwxyvPpfiVo0JWGbot16M5HuT0fsnvjjOPtF9X5OyX
Pej5NhiXpFNWsogo9yYL/uewpFjS2NP+/JXUu+vJ1EKC2KTPU1ZKyYm73WQ/nGq0RNq94Y2kP4BQ
bAhFiXq3Txux7ggF3NUg8bOPu2kn853pUwlpBT1yO05QeGBda4j9mj8c6UtA/Pmm2Oh8I/k+1pdn
n3ZyzUy57lMPHOkNlZla7sMMgIGrUq6uZkq33kOcxx/40lydxHzmbZjp0weh/jcPsbP0/t4XkAuA
Ox96auZxp/Bh/4gzVDlOIdzoDvlFzJs62zdxmIoZkMlijOvZ50Uh1ed4irHPJiGFXNZRtWwiPues
A59jBNfIgUoF4ghCCgvAAr2HnMmBtz9+gBKknBXNZG3z2qLcfRoSYSXlw+xXbkS6dJ08mVsi8YYi
kt6BGyNOn56JD0WvVj9WSg2lWTZu+QSUtPqR2PV8RscYIT98Zt4W3b2fbF2aB/SLNwkEvs7aL7ku
kY7J0c8HOZ5+W3sLUwJT/LJmZBgYvyK0bS1Y3ld9c/3v2NvbwmwIMQlJeJPvh5QzXx3wTsBEoRoy
2M9VPdhecis1Q5sY6m+WviQN09pbanqLhBo46GQzKOSOwyCzUYWgVVE2Z9pxUAMnUdrsY9mzTDfz
JYUxPV+gZLeKonYTGX/gxissLxz5H3yVrS7TXanD+ZXxcErqydhvGszQYpenFB25IsZShGhIjp98
cWYPx1P6vVqiiN5rdqH8i5SxBGtbgr3SdFuvHXBRXvr65stc9DPvNLiBg4xSr8sKgi3ajRuI6Vmg
cfEEkOqov0VI4Q3nALR/QMealuny2lqoElRhrfBxrmKhYQ9ZE5+RrYznP25EbHGHd3S7bNaiU6TO
7sQ9JTdER4XKa2rpTe5fJYF3DCZl80088Wds9c73YBz+XP728+0vkX0dRx+S8O7+MwD1ZVU0aCDA
KmXaBWlLzOkKrnL14gwJXDcp9wriOBnV1hs7YDIW4r/aNgWgiDLMPbxuPXLUSGWYlZyMEzdyqsWk
20TXYslaQpQyrXIJlaIFaPrzH57mLxS08c7+rK7x4YwK9cZx1OjV3ncI+1wPz0q9YTvzAR/FsusK
4QBGMnX6FYVlwDzLc5PQRTWOnQRR/DcUe+eN0Ht7zOBqhF+BRmy6M8LX6sNHRUfHWQO3whEJdchv
AnPFaz6UNqx2Ls1CAQ78gRWAeGyeMY8cKgAvuUQCEpNUidyp4I7EUo74/xZCMg1nJFkDeS2xEBme
llinR3Gozr1s5I52/2f8wf19BCfyFzHvhiqZ/H3A4GfQ2rTUFRSYqBpcJembV0T6eah+L7Fs50aM
MUTqw8bnIW0LNrBlBnjoGqoGEy2moAUt+cuBhi9bNKk7qa/+6cG3PBSEouCAZVleYQd9DgecB9Sg
ni32PspR2ZlOtMEw0aXAD8JO1ags0o1IfiQfmDPWf6i0QgYTgSGjR16RjOf5SWf/fniuzioUlcaK
Si9Y4+zprrJn/EipTonA/YNhtwqis+lUCKOA0wArK8rs8kCcCDzEHk2ozLMx2uGnkflxPwBuOBTd
2sW+znJEuwvVEW3wTqtzpnZvlyBFDJZ85cHt9q8Sxu4UGtECDGBtfkmCKYPoQU+F+oVES/HWNZfW
kFD8G0LIeqK6XqCYJW2DSj2ptMOxDKMiP+fn8jxfOAtxxm/DFZkUD2hxn3ifZraz3iwBq4liAj+k
jL330fBREYVsrpYOUVrEDzqm7zoAXdzyqYR0iu2YG4Ysoee/cNL6CYJ5z25ObV/x0K/pAbriKHDG
Pqni+jtAtcirrFVRM2Zq6GMqt94DV7V+w7UilCqaGW2J+qAbb/CDU0mkPWgyRoMaCLdERgxICTQi
olTlGcokIAIIz1HiNQ6Z7d2LtOgPH/E+Y7bxAosAnViW0NW8AAx8+zTWZQvVVFpgLOuWO+znVk2l
Ml1wGjq5M4hhy5OvOiMvIadl346aCy61v2uMuaLDsHIX5lvIYvit/Hq5kg7fYl/rXHzXdPs62788
+kU3V/0+1Ugo9rMp3hJ/z+ET5mmuDyk5KaikeJrtDEJpNVR2Z9tsrSd09jx70TA1vwacOXWZuzdR
SOaD5m7eGAAb+3TAXIE5ipc1Dd2E8OkBKTl3LV4fiQ64FZjf8qAjCVGOe+4z+v3lJFrfH5i1slNg
co80M5Sgm8FOcBltaFJKOhhdXfmIBplpBaxsHkRs/tZ1lM6u8K0ogPN1HG+kQEkLQYp34y/W67gv
qJwmsajK/i0RQFfi1svFxOFcxIvVutbCwbvFlLcNqQlhuKguveVNqniSAOUfaBE2OkTrUPnJXa7h
HMMCLPNL58vgxeCgAJIhHUsYCBw21iZ9Jvs/PLNyhJf0C+qoXaA1GgIou2jLT31kxnR8M2L238p7
/e2H/wboklrsnkAlv4GwTb8Ed1m9raOAozDea3eDvjE5YOR2ev2b0v61Mj4MtKeb7+wtKWcy58Tr
uqyINPuZCagWpIdaI/utcwpSj3VKVhxeUmW/sRZbbMCSnkDcPxqZrvGNGNomwtC/PZ8/DmsqvLZk
/kyhR0HlAk3uo578lblsrHLvlchKHNgMy8Jm/q40ZNs5mpZYxQiBAxXeizrUia3nYt27n+Uugklj
nbeVFsxcy95yhUz8oD8AJp5INMMKqzAS25QzHuSpc44s2OlVBnioxFCJEgSPQyeJaxkLzLRjlmqv
2w2doyBlrrU1Dk3yLsGRRsDaob+9twpfJbO5AxgLlIRhtiTWGADHw0Be5jLf2dE6B+pUcfjZPenK
E/rA5/LUX/C72e6q3LsxI3XsBd49vFdYjIMa6NYf0zwlfL6BaGLbBo8WFppmOZZB/zgdw18mVgZR
pnnXi3IjegBfVhDHpaTcEhCfjL+sN0FNqNiYFLUAGFQg/eL3udmJLQlyRFWcJjlRPPzpstZKN6gn
u5dGYJhrZKfPJnzn4oqHYsFJafvtyDAJm9UKehdzmL3ucv65/Ylac8mzpnhQ9RMhZmn7JPfgk7W0
kGclckdI6rQpsZ8StZE72vDTHj726yIL+91gdBEhPibGcX1Xva7nNNe2Ydso0XAMoE9eNDFqi7gI
BEA7/OJIJRZwP+Ij6zLrexLTbN7T2chXLuIexs4SY9//OoYimkQb900kzyECNnBVjFDIUC8BegI6
meF1FWZ68lbzL+spFDo639PjcV1U3rWrbcNpEEa3td/Q+9ZmHwF31Z7brApKMQ/hU5EOBu3O7cP1
tyc72XsHwL6btomAZtzdw+TzbU9VroPHWwO1mJt6faY6Z7vrSNVCVMs7EiOiOup9Oav+B3lx+ED2
wAD51ia2uUh9Q+wSPO30zmkEc28WlkF13qhLp5Aj1W06om5OFpZnHyU+R0rrIhFcFwxrQum2l0L0
FPd7zOmZF6z3iycwmWXxUk6upyYB6JGERSiMXxqmz8uPuZ7/V9HDOtsv9MS2C81C6stRcvWxoMPF
Rn5xJdSMYpsKr/pvOsNeMpPc0rVqox1DC8TQ3tUIyoa+wTCGhlU4+IicpPlFK76wqaivIjoI3imf
ZUVyHePHp8BTbr90uK45Nh2xc3gwbbiTEM6VfpP8OUQ0n3Imyv7vT8roUhYy8HBq/bi0PDcRtHNg
yX9HXZSmoTjbFYom01wmUQt9zDVRUvuixzvqvQA2PfHWnJqHg5+CoXcLlgxxkegOx0wafgkG3CHf
ZcJ3sYeTyR3Wrpkew+f4VM0DPwReXNhw2G/alKaovttQ1pUe7G1yLrMQ7R7qn+c+oW2n3JlT5Fg3
Zkb3/kUTnpX8Wl7R1C06o00Js+t2ZzDGxjNiAo7d2FhtSh53I22DWJMtQ+pw3Fy0rYRxq+aiTxHy
h0pap599g2q12+My93UF6UC3cIJWCEz22NNDHlbg0SJxfxptYWpN4AQXL/Z83Mkhl0EVq8iMTpMj
S3ytH7B4mpL329YJHDehbGQUTD5kWU1cOl6XMtFDN7aR3jhphp0pYc5ICsI+gsFbLbnhdC30WSLs
Yec3LxOgDoct5Z7dKCasWktUnqYdDahaJEJkp2jvMmjX2tlYBsxO21d4QkNWDqRFY+bj7E5mE2nD
S2rPAmc6N+39XHoYPl27eJcBbJwv3q6X5CTdTMCB6PGQwjVzI/Qwacjc0m4tHI5jPlJengtY3Nsp
QZRaBEqnhO0PVAXpEdx71gWF9IGn5LYYc3TwQBfJ4y3nOZAsxFJeNx75DjUXoBNePpNq3wJs1ZYZ
GzyDxj6+KCIAW+eOn7IQqGuvN159giRlqsBDKiLUl/iNvOiGNCKWIWQ2LFB5teNz4Z7OkhVWW9i/
PUTzgniCpK65t1QqtGsyIqQiruolV0h9UiHiShzUJiuGEGeK8Ah+hxBrHXRXljUdHT4VKQkOzHuc
gIDBoPKQZYdCrEHbFo4O9PFKN+b2YMim20Bs165REFpCQ00goCY1lrW1iQgmE8nujyJUMDriBXMT
vjM3DEVPp94GkFh/mnl2fH0jqAJNiygG0sNgKQGLyB3Wa6LxapFgLMCIvcuvN4LUy79fgGlxuaI/
dUSr5+B/OwFdgjVjDx1dRPXnvXWpwvA83hmxAdq08oPXQJ9iCpLaTuhDZvz/7OJ09/i8EiCFN2Tf
z+4RK4VUHSEChtbme+QBrxJc922rybKB+4FPNP0G5zr8oOTvBaYDT/KqTPlno2tONNEGysfO2mgJ
tzZcCIPdISrPy+6JF7ZTWzaN9ozh2qyKk68vjzFOBDUVO4149PAOQwmcuilyuFwRmPA+ASv5rIE3
UZ0689zZuN0SQztJJNOrTYZNzOdxsEBda7c6ddpGC3cHKfrCJqXRIpAA/E1o1nm+r+fffacDRBM7
kFApmiDaCMTRuK9KmaSXBksw7H7m7vBjlXxtP2LgNM4rGzOxzwrNlWav3JXOHwz1N/Svl/EdsXPa
VM8SoWFB8h6/bchZ24NvX0fHbxdgkJdZgLzZecvgmLV7FWWLDoONWMzrDge41PV6M4T5bOq7WsAg
uzSDGYe7lMH15vzQ2rwiETEjU8MSMSrvztVkoQmmGdnR5HIaF7YvzbUvB/vWU2yHMBCmko9C1Zzk
gy0+Y0yfEuUhHKzXkyBEdtMYwKatsObkEbdsrx9zLYClAt+ImslahHbMKq5Ps4AX4HKd6JY3txTv
kL5Yh1aF3KqcnuZXEzC8n/oAEXDj+oe19WWdjnagmHBuJe1M0De+gc4gX+g/texSqGHa9tMq4y/z
PmyxuxQ99EFcAdFl9Szn1boCjD9oBORQ1W8WHdBYW8nyQyqEfzEcHaqk2y4WhPahzF3FZWslksgH
3Yc315Ns79SwrrVJaRC1/I5S5GdgJMg3LQAKOkVY2ob57Arz2JWJC7vCRBJr//PmsyFt3zxRVMKP
KNzDRVGo9z3DELcR1SvNO738V+WdbLpejv5QHYx5mr2A/4q1BH9eLrAA3sQvxlIZHQvi4Nf7uOGC
by74bH4iTF8LJ7dW39S5l2fDiEy2npjtdmUxIxPtFD2IqTFfnYFTUOCuJQtZ8ncyUwCRMSXILHIW
JdM29xhf6dbaDqDfVZVI4nX32nvVIjm/7h4tAya0wGt1BlXampITTB29fE5ZJL26/Y6MybFBYLzz
T4pjNY+Z3tQMBn2gPxCFV9nkUeKMftOMrSkVDsPi1eM2pBzb+iWggwNG0R4v7ZL/Us4z3DqnQGyz
9cYm5e/OJdYz8wlgCMsfNAj84M8JCc8s+IL1uoMlpF5oJgEFwpgx3ekiMxqXyAZhgD4USRwyikML
Db1vc6db9QsCe3fW+JxPfDw96zZ5XblZe/KDyzz+gRCE6UwtrFbeAcHV//0yF3ssMP/jMbHFU1yC
4xfX826ed1m03ySqQbEHtBa29h1DVMVu6JbTm4eJjluhUUWaElgIsyrVVIRBp+1iD9vp8qMtsuqi
ogDOX+e5Zpolh66ygVliOZDHrRzMY4aVMeIhmfDaiJSCmCtL8p3w066pakMf506QK3aDHejtv/Bt
eOX2KkD0XEM65zSQn20R6p1SDLAfZ6fZhNhYPof4Mx+Jn9MlUe3PgU9J9Fb4UZcSObF8bw3UhyIs
GWlvI+R2sEUk4HvE+9Co1D9X2gpkKh4S5RJPy94n8pj1gcJiL4hEMTucjo40xRDZQg93I3vK/2ju
5XCnH0vHcfkfs9buILwv/0TFhvKVSNjBk7J+m1slEp075FsWuMOmQH8ML7OKGFv9Q+TNceQA8g87
6tvC8wn4ispQUbh8+ZZsPHkbv2p7HjiRPfhLA3LLQX9sJnihFQ/BQeXy4BoAhD+JP60iHTRVeR+I
h9Pi4HQ5gClrSD+MnjzPCORi4Ix90rHgT1+nGMwzCXYwY7rD6Jm1LcfJ9qNv0B7Bt4UhAy0lRJYd
/mY1Y6w4DqDFGK7K4hTHSa9EgrcwRjCytZ6HkEVyFAol0e9QGRAsWYrup7sibMVI4Oh/sO6HoVNQ
TXmBBQ4Ni3tmeLuH4HtVxeiHrcZXVwrPuwAmuogBKm4ojlPw56+BlnqBt/hlJcZQ3jL+y7nWrC3r
HrPm1+9OoktjWCNX2ypXK9nmJNOWxI3JJ0psRrmwYgesPyUoZwyIe+rM+8Qj3/Lr3GFxYZr+2ASH
X0XDkKD6HAHs+ua6dacCFHLkUXiP7b1Z0hJoau5+KtuUCApuAUpqJZO7OW/iE1rY6GSEYtnvCpjz
PKsb+6Op1nQW6UI6Pl3ZXuvqVyWvHJ3YMPHo0vtTV7WUMb98VwQi5kyWGtdcm+1n/FaQ3b5hiIf9
Vik2Ik04tV1vwkhORY2if6x94SGGdfrnPphxGNWctOdBZ8y5oZnHRYcHlN/9liqZPwYFQC9oZ826
wyRc7A1lX2nhVh55rrCTW030MmWMR8tOI9TKEgTjtscQFqrYj93B5zPOq8z0eIB92X0D+xqj3caO
Ga4a6NCmUdusqIuglpSk4c/X9AuF4i5iQCRVthHE/o1hbEwru7iKAbpX5a8TD1FSLxRrYZAHGVq8
LRzCDy12PjUokQbAq7VlJMGfD9B1riU/+qxJUb4A6LAHKwLE8ddIsT6zMDzdkqYZn+UP74KUQ5hw
e2bIBjspLItLhNymIt84nSlB0qL9d+ZP+l9BkBMjq28+JzhjgPlz+QxeTlnluF9MDPUKGBCdM3oQ
kNIG/i9SyGcqRF03tU72EKsXO9nLn5DxhdPB/F5JAuGvRNdAUdgkKpz065Jcr5fY2u7MfKNzK5OB
alS2XuaAJw++JEJr1QsulyccHwIcMWRgOrtPbpgLfyiL7HNXOw2LtaP0nhUPjIpK+pLl+HkdEUCf
FrrugKnMD6WII8PNqhswaQW8BGEjcaTTro7FWkZRYxUfyofcDSgESfhM/zg0X9o3nbRGMiBxCjoY
FYBtP4q4dbfJR2eAPqlr2vURO3buPs2oXv+WdfwhQNHxhWTe5iaIt4yE7m1DMBD134BTS/R8PuA/
JL8tgk48XXj3H2PmhWBHEBeAwJTs9KyfKk5ni/BDvKK3I1HjhFzgVho/P8D4Jhk/xWr7cvlsK3Bg
vwF9SKCb/5zq84LALQYU9iItJL014ReHavPH9W0vlNBuxl7Glu2MBJze39KwNyEGWsNXEx5ihpNV
LXu1xKMB/RQxdg2nqX8a7OsgOdX93x9eBqqPA/Ft1L4lr2cgGQPkxKOm9jLDVykWfyli37l2tdss
nt9hgLkDm0nSCuAQWbRcYAk9VH2y6+HRCbpk1HkPU0YZQdk1z4mNVUdAvQXMa5aGsSnVcLkITwVr
JfFQTBUqdCxG5j6pVWlHlc2c+Q14mkiy9WwWAbcBow06brtmkU7p2VczdwLI7riwMYnBW+XGal74
98R6QEwi4DDfV21LDkzUvCAQOcep9sRRO0AaKwI2Q2d4uaYJCZR6Xn/TsPtMcZTpx8qUJOE42I/m
Xzdl0E2jWdC8GQe6++QDgLEfhl+StTNvEHBwup15OCv2O1yyLb0Vbiz+/fqk0UDeOdDOxhDZUI3+
ejo2uwbBaBC6jyMw/CKVNr6PxK05sBmrzRXWPBjoZtI2bBXNnY7RAd2zrRlw9+2baahIZ+wYyO45
fK7Y6DCKsKwbNmxurJBw9h21brCVF65+xkZGLXj4GBFug3HsiOIMei3HSYcGdPd9q3aA2iuZ8DEe
BCdn2OOeDHE46jdcXj1yBnjBSw18Em6YtiOZjEXLXeJbXQSHrNaPR48979kZRDKRs4eyBgaiVFqy
2kpqMLPbS4oj4RWKX/y5ofTG+P+hMpR3opBOwuNBQC8iSEtSmZjC7hZFaAQtHVNMOKhpjXPmjCtX
/0/Ww4A0HWeBcGN9OPQaf6aHGosU/FbO03FQbVkw0Set2YDIinj6wl3TBAwf6yWJz3qdqwWMHDyk
9q5rxKdGWA3Qs4a3I1adbKodv0GefIFXWhgLO2QavfuiDdna8j0RksmwVBRNQYvbBXsvEcToxXjC
7N/t0qYS4x3JZGTrZWkl14W/Xa1NE33AJQz2rrP+msr9IZy8mpf39B4qU73ok4bNEOEw3N7nbPfT
fn965OiDCbJ9WhZaOviF1XFbnIO0j0QZ37d+T2A+FlAnZ1cFBPyEoB6SiYEDSd3dQfEChF986B/p
yr5s4K+rsK9McqfQNO1QlnT9gIzG9LVwrP5JEI+HGYW4GKts13eoxmtJEgwq8kFyFkyRgifnVKj0
mjCJypeMip1TV+4Me6EgoqhBV9GPCfPKbJ4AKpSTbhAcrRytwY0enugvjGtM1eB2LGtTuzk56UwV
zsNyBsS8IzsOdvNxcjIgOT/JlAI9btlW8ncoTAzFNhh4gmoMTTZc67NPDvIH79dUSwPc1ie3VMMp
dsiX4D0Jv0LztvyzVJodPBnmD6DvPSSJqaChIrvtFBC+dx+3DTLI/WJqhekhC1MeqIWHcOPMOXOO
rF+Zc/XkvSbyg2XTToOxBZPfG0H4wfmhxWU/WfbqzsDp0H70gdHrTE7IePBF6vQ3h0KCtdqPFnAY
E88Rx1ZBirGRAtFrrH78ca887MENdE7LwnEej10dgrmAsBJpVgIlQncdz0bl8CSBz/xVpmmwgsDC
n5dgHy7clG530w796s/70DI/I3JRrbrTFb5KS29ruJjUEV6VwMwva/ongDgZLVjPayYI5pdnk2IT
eZVn+SrILozXJPvzIDZaNIKSte8WEQ+5XvqDgG7Y/1fvW95NqGIjFp4Y/e0lZQCohT632u1mDyqY
M2c7gJtEaMSiDGN9wuZ/OIl4u654UESaQnNbRlRApbbKCRyd2EITDcn+phY5P/A5J04Ij3ukmGVY
/5zB3ZvPAmJfZHNaArH00r5XtIGu2Z+lGcoXc/rK4Qw5Je9YgBSslLO6FRZ2+LtkaiJ3SbD+8bSA
Hi8AHsG6nasUmgX2oqGjpbLq8q9CDQMP4rdlOCaXlSKt4KW2AK3HykRykvC/vxmaLqFucCt8WA2m
wYcSWLP1bXwb2VrvVixveIqhlVdyan59I+LXdtvVM+/fjtnaswTwYJuvimEHv6CdCjfIbfn95RyP
t+jsXogH2bc0qRocj5FizwPehFGzyn9uRP60TT6YyAThRZ0yua9bLgY7m9GLP+WeZwph+XRXWq46
y7BLcfDIbOW5B26Hi+Z+m9rIMcDyIk383iRJ123wOo0ZNQvAH+EP5mmiqQ1U8d6GXVlI2BvOJcdg
yFa6wCrKibzuYH964n4zesImidTF8PKZUaY9hulCCHSGvQp7fRuVYz80Ca92zUB1JDXvv4dDXs4f
+DaiPYxKgmqrNGN+ktySye7S2h/T3gPvOGYxtAHBfjhGjwLuj/qzYhHjFaxPtOEVuwlUS8W078M6
/WGJ1k7GF2cmMrmN5LNZnVqKUIdJ0XtmaV2x8n/pY+t3qjoHCSsGIuOzIz96BA9c/zgxR5gPidMz
5xvaCj117ec2cqunuDjF8uKnRe6F2CP7RF8xBnQzI0VHTO/O9JvTX2j/TAM8VhbUthwegJGJfhtG
XM9HpL44NJCLuR3o3VjfVGHuk5Dvlh6zzms8N+gar1JH0bx+AOtZMhmqoef+H7YMzO5kDjStnjHb
PW8x8iXQbqsXnQFaLEjuAfU8y18mFSd8SHjfyM1mbYkQcM6zShTN/RXWaMjhR8KMs2gyNhxQq019
Jwm+awsabK7rM0paNwo3T66IthEtzx6RCPxVdLWjlPwT1i2TQF/ebN4B+xhQjqBbv6898QY8nvVB
EVR711wBpjwsuEGLW9UulYZG1ehrr6JwzGJNvmvfyvG8lZKJ13vjRcqPPBr4YqhbMODkEruJ9lZx
5/GO0G8JvbrpGNuaRIDSRPjvn4P22OhNe+7qP3DlZZ7ipurhyo0zAcZmM7JmWI4/htQMwyaiEZaa
i9CfZ0W/KajCZS5Q5F41m0M2vT8/TMtqhn8d5WQtVCBHU850gGsI+A6ylj/l/Qx5flfcHmXbJy17
HeZLEkL+hT08CEnEkLltjej6sVbOhbK7XCt6nnhu6itko8n8jTE4WZ1mfs3cSooEXC67f5Fv2IRn
BdrvgsVOAuIaIGJgU3yV30CqUrDBFXLVPddzlXqPmOTCNIfRyIoTb91w5j0UovcEfB/fIQlXgiLN
6KIcgrzoBVbFAMgPThi82LAmChCxHSW6Rdte6aS2iaJ8dkcQku9008YjOCKmOLhs3Tjybhz5ImUG
iOsKn4C4e/DfKwNHw/pUMXB+qms7nVbfZbJXxaa7S5LZE6shV79oIRAr2ATVGJOVTqWxFXyw9NcV
fPGLChPaflDDw3Ukr++zcRJWGQa9DvRej4hlL38gpjf5Vdi/78xHV5yL/h948Hc59MY1UbVl3VUB
OOaVkIM0j6r8t+9PDu27j37Pqj08uVg9h5uto2C3yiLmSX3PPxA8j0MTui2IjtCJ15Nj4OrXgRQs
1/dLGfhf6vpGd2aGOTy5GFV3rOIz9cgFd49oobwq8bdYRTSlYX+CTxXBk+XkD+Fs30V7aqd3LsOh
G83uRPDuQePly45yXXDqmnhAEzJvZnCxOGdMufc5yBH1jt1HrFW10V4R0UkAKGwQVSSvDGtltWas
YLcwMk6IHRiV6Cr2DCIDnP5xOYomj6AkhrQ9x9+yoUAgOXjXdUe60jlyh7d7rah2SAnMNvwNOQ64
PT1JLKYSkzPoKwa0MfCkmPeTaX4jnRz8QBb3OkYq3vMzLG4GaHQWiIl0DOpzLbSA01DQejTjpBD1
8KG8eMZxum9Jr6ZnOnuzI537rxTLTiWDQsTWJoQFK5JVaPffJVT1+z4WLCHimx00/5rhVlJum+gN
51kPimQuoLI23qn/Xw82AsHaIzikLdczzz68WdcTH2SpyqbklNRY4D9n5xrH2XymldzB+Tjo5aJ/
kUvaYbF8YPyI6utkT95LrbTG9Zq32GlT1dnIy8yLxWUMSo9GtP8b+KCMPJ8gkPUT+4GnVkmzjW38
s+vHUmu5kqEDH4QBwkSBM6t4ZkVA0hRuOvBB5lqeS0XzsSVcl3CJAtKnmYIrVEdW9vBU2Zio97Qj
7kb0JrqQzeN1pLZSsk32x813J6uyrpP41HyYrLD2uJXE1xuwFP8tG16GiOklcQ7Q2KR0K+M0soJH
BDGwfDHizOOKnoPUu6JJXkvCcTM8jll+u7LEqeDwrBNtLA3xX2Fr2ePpwy/Gmthqhd/PlNO3oq8p
PvOncjiD0o20+XwUegPv0TZVxicRoIS7rNKMJORvqAaLF4e6pna3Osrf4GKW/2imL8VnC8lFA+VR
ZMll5tVp2hmQM/Ov8vZwk0eFP+PnXRpjrYAnWxEIPkaW/LxyfmIKevcLX+Ax0WXPJ/kbYTexCquD
hQpJVnxEOZrWW3uNsX6+GjtU3/5TBi2DUvhMVzp0IEREZH9GCDuoyWklGSEt973GuszMgvTWSdDP
x1nYxrlmnJ33ov9IUNMB73V2HOsKrV/uNigxHH2M7z4ePxRBJhQ3Ra4HtnGL7gTl/09G9KSCI+o2
diRSjAqmyxgek+gQJgiT+9ltTTfxHTMDoW3FCSQKsbAPrfFpueJmh15kJ/otyllUEsV9lEdu8RJM
LAX/c2OxHgXW5Z5VRcVKHgxYJc+jg1HSB5K5FJaZBmhJr9rLdYYAxQ4vRy3OyPuSt0h2SdJyVeef
tgOqCZaGS7qqPzQBKpETTXFvW0igf6fThc45TaRmMOsNcgpNqAeBNtXk2BfjiYbLz2FIyPu0hPkG
EB8E1pNtOH06WeFrKfh5WcOJ1SOtSypCIOt5HfRo0Eifk2s5GmpRyxOpIPd8xg420nMdvT7HJihn
SACSaHEBqURQVW7XYP5nu0cizcXxiqC/n/HlU03VwZrbECoYsowTsIUid1RgS63yZmVfHRzwIUhb
LhA8bM8eBrc5IfVgTVvCH/sXEOJnxPbuDXmIlO8vtusJVwMJMKPAZHWr3S2P/cCmc8VKjlyVLNqn
0IoRZxVIZwTS/g4mOEuJpayPD7oG2lgRtrtRwvN84JyJjtIjz06MXiuG0Ip64CZQ+B0ZCwdSjdU7
+ifror/noklJOr9Rkla28GKu9CPKK4JvBm7oAF9lRjLBdUcqtwkguFV8cK2F8xz08VDQgRxDR0yr
pSel9b2pVj3srxWgK1bq28sSvX1iNza6+iJGpCN2HEB1FF9CcKA0NYC7e/Qm7jUH3fCB3Annfi72
NP+s2iJ9m/k1LUOh2EihOLUVCWNK1MC935Zvvw3s4HFEHdkcB6ubjzJG0eUoJFuEqk5eDYG1/X30
3T35XyZIdailuPXXWErJ2DLOCabNv1++6VUKdF+OD1NQ3lXxvzyX3VXjr2apA9mVT4aTg7ltDC3j
43YLz/dP/ANSZSobXeg8bg+bPVF6GNXPi/Ov5zMK+DK479SKGScxS1aevONX0ZICn641zPryS5HC
hedhAJbJTJU53XcMxJnmxOX5y3VQnZNzI8bn5EWLtAr75UZZ9JHUMd4xJ1rvSxsevlRDqi7SLXDw
0tb7FpjNe9Nl5dCZTPl9aD2+tmbWgp6pld0oCprmEsbKbxzITEZ+KVvryY70lokEQmg61TtGJoUt
gIRzxuaIJCK7OSfY8HOo9BeTJMAE+2jBqvetxctvEc+akj7e7L43We0PScreR9y13tTxLqKZ0HwD
OsZJqjXtfpxSe1Lcfdq5aQNipBWPahBcSErIhXnKbpH72YLVpzsBexQeA0DcAvplJwTUyz/9t3FH
Rq51LQpYrVEbZwriSWMNtKU6Ds7B2ZdL9APGtK7fq0ybM8QOPZKtoiW2l0wepsIAfcyxFgHLxYYy
iFywFe2aDxB1lPWoHkoA75mwdGZKcvGWc2OCukH61beIFEJTGpy3Nqc9Ktr5Ar+UbLiD4n6gDMz3
+9sK17V3brrCPKsyB1g8jZcVt6GE6f8Wu6xwSVO+Yh8NOx5Q/jcC/mIiYJ6UXGFc5LXRMHDtqfxG
jQ1zr65cUkg5y/ssk4hF5sAkVqYXi3nWhrFphR1v+HwJH/N46h5XI/Qd665N9lglNVXexGc2RuaP
+ZNGtFcB968CeLv189KPm0sZSL/Yy4V0gFkyxH0IaqG6VniiHpUc5vQJWJ8AjJMNP7htdBrPaHDl
st50GvDBKa6zkD7KD9xCtSyVeyORTThDu3eT1gY2dg7om4g1sUlxSzmJiuhzhxn/3ZpbfcR+F/aE
vTcVQOyjToIYjJAhd0MZjxUQKgl774R3tS9tp2U4RyzVejv0vczmaUFlyvpJ5phB+3LMVwlXy2C3
Zs69VtXiEk75Zj2rdtxqBRdjyeL+xtsVcASnpIcvf4ys/7ubD42GBulSozirDAMXdzTdYnYcNG88
PdWFvN1GA6zF2KDshOcBAzV2V7suChk4Q8FYjErwMLG+b8onFuWOJuAlCeHYprERVqBWXEmuXyRx
BXAS6AgugwilJWW4QLlQ9SI9eDDi/oe+L/TI40m4uT7FxqDZi5kaXZ5dm6ElCiRA/DrICIW8i3g7
FQx7RHpjb2MaKJVOvQzW+bxFmXIgEu/xnoOpxDp8Etqxf14jK0Aw58ZkrXIQeDjNcsejNLnzyBY2
5knxO7bYqiO4vm9782MZ5NyN03/R1559LExJrTZbSAiatupHwykNCC/sNLJtZxM2U/sq/s4Q8ay6
0xKFSmNr1DlqqJm6nrc03hoMzd6fO6g/ulbkdq8F15HxLNWyWy+KWm1B3ZDdctMOOSTxvljrP7OB
BnP/QA+V/QBj0zYDlq2mS3Ocr8OjlHrquzT/c9mHRDdH1GkvGeWohocJgpuBhnDUOB6hM/RbKRBG
O4uY2YNgeE+g8993ad+/zWWovEa9IZqvqRzurF7yc5DSMxR8FIe2cSjYkZjN1gUH5R4uts2u7nO1
EB1pCsQNzMPPWBbPeqgXh9F0F7SXYL3Z6fxQxCV0zERqeYDjt6X62D4hmqTw0OPLVHBKHqKMAtcL
6I+sm4lx1t8z3UvG/eVZiDOCb9A9YxTarljCl0WIfcpzT9K7IYwrAI+QK7uZV6iWXntSYX+SoZ2F
QeWKJ4yhucn/vGYml1ECl5gqEeNY1pbVnfNNizds74xjz7ijfWCcXsoyQwNTJrNvQS+6qgq4xqO6
72SzAdb/Tn6j5m6Kkv0c+yPoNNLhU0Llsah0MkJChPwmQToJnHNjSDgsvnKdMgwEe1ifl1i0mNKZ
Mhv1zBo+vE8LguMkT4ePG/CZMZhqR55qcRNo82ORfPgJUbXfiOsDk4Ff5JBwGbDjA3B43E3PeXpK
qBJe18WtVovnbj1EBdSSds7ZisRVolMgSYllZL2G1SuwVOGzJt7kGyP5gFJ7LOE/+DjEJTcX7IO0
C7yxfatbNRpaJSliwP3ojz43UZbkFS9YT+M56SRaZQUlQ6fYlXGM9izMaHcUdajMMSmcShumqjpc
HyZmD2qvQtnC9pJ4Mtmg5cIHphNrSnvhwq5G87TeMDASXWx3XHXv2R+XSl0ysFWEtPHq3MbU+w0D
lDd9VkrmqD6e1gd7jCdIvvd5DRqlfdkqr25siz5KlslvN0oQxNKmTD/GRTtE5v8ymdeXrxiDO3Dy
ApLtykjPrE1ywGRQPJBkLE/xuLuqsHhtkl5MKF/HtbW2JMcqDSRIMnFzP/1KusTzgpd92WW/YEmn
eCCbXoWTPa+Upqyd91SzzKjoHE7tpu1cfV2j1NmNhip9fsFzt55Xtj0K/ANv5Go/qrnmKGVNAcaH
FJMwtwsNusCgmIya9LN/5Npiur3tfKN37LP3dhST+QmP8OLuH7hwMVAXcddT3DLG4kf2k2l7HRW7
7sI7dRzD35JMQvyw4K5F7K1tnvCBJkyhRgXZXhDp6JpG3l78u00XwY2j1vkUVHaWIsAl7V6Ga5RH
vAN6zJRP6A4JjzdBakigi9LLfYStka/DzKC/6X9vvzVr6JP1xB54dYaPHOoWbTv+ME5shHVhRaY8
VfLeUuI/8VJKHewR2KPslPlpnscrFL6CbaSXhL8JFx8E8Fz5JvShUJZbaI4QBpKQkXtWCortJwx3
NXpVX7hJ83XXK1FGcUTx+njbH08/nRedHqFx4FzIokd/PH6jSWnleutmSZrWebOtwm5ZaNM8maoK
2J8jdpTFHJZi0umXOXmgLVysHf96wKtvrUL062ONeABCbYRCBJXEbBoE+GRCr22qUyW+LLUUYH6T
iJpQk2UGEbKfnzXtjOBi8n02N17DmRtukMhsuDbxHQ//NrmXlw/kOsl8R+pl+Qhbuo7QMABXwpqP
EKp/KJamSny03j5pGmRrsoNM/83eNm288srUe9uUC4nsOFL9TKNVCSbmxvpgSpt/AVXQ81JtyVaR
MXUJDeBAm68/pYoY5mUmSR9yD0//Io4hm8OCcD7oT5rVGNWJppKxX0n+bJZ0M18rOlKrVGT37qUj
a6umzE4kJUpOOLxRQq9cIqx26MmKrD5t+6dClH0nspPHAl4gArCoSyFDYdtAJGGN2d15jHNeR5ji
RjPFrjQ4IBFauDlppISEZuuCgXOn7rs/Hjy+gdOApCjCrMVgnBKJuDWhdB+IJzeyQ/yQhhO6Vt/D
XYqeFq5LEAE+nChEFLwNBJHOMeNHSlBJSRzA+chAdjXnjKHA0kn2Qo2g+V2M2tgKWFi89NJKGUD/
EK9DUHN4oksglHfcpOhfJQHtmiz/edLGLMU81L1oDC5xORLjp+MwYJgIMjrEEAThTyCnn99O6lGK
349Bn6gf2+k06n/hy7Pll3iAr1o8Aq8P9YVxnwTRs5NpjfuafnIgsMFYeEG58tVklxEz3M8nmuXV
mIo4y0kPmaW7nbVSja1gNXYyn2wRi8C/8zMP18Us5cXbh3syzVPzpxoZ26TPKuDsxdsXGHt9tCM/
Nobx6F0TtwBYqn5Pr9zysjcQZSfFIMSpVIXVEfWTKsMhJeinPRkegu491wQs/HNcu3GYvBnCVPi/
sK3TIGVgxdkWfXkRrMqmByRP7RQpf28TXcLObqxnKuuQkbWbmbT6FRt6Lq6UDl/hX6Nn/cdGWfek
a6hLQebimwOsY3VLr5IJ0FatryjD1ChOrf6SYRvDeI6P4ZQ7dVPF57x8wdprVBiIAkFw1y31zEw2
YO3PizAa6yCjQ+zmjCb+OxOdDtXaRPmzMlCcMdMhliTRau24dOoiu33AovUGerV0oJKLeUCHTsnY
JN4vWiUPLOr1LAQhwQehK9Z+8S01R9cQi1LA7pSN4DiqbmlIgdTBWYlB7Dvau2B4Qqx1A0+p+53s
2kPTxT/uCC4hBIl4VbS0jYffvTBYXPJxjHmtZ4KBCHJT/p5CF2wz/daIKoE8MNhMeAtqawRbjOn7
hR1AYrHYeNJqsqJW/jc9pk7KfCj3bAM0YGmEDwLH7vNni5D1/I7CuwV6OoKD3S/NprgzihBIEuSX
PPbtlP77mlB1rfgBX5FRmdY6bDA1BMyqJh0WU5ecCirbHOnRWd9a+vlqS+F/zD2i5j9E3ZDe7fZi
RrUiLXq4yPSZ/SIsqeXu01bGIYGmOJOhulQ9ELcEYK52JG8gZp58vzo5MOUX15n4/Rbf+QTglcm/
czaOgu2nk4kfYAMBCmJP6vbJWOLS0+cXRpjwGhzL03eeEV9nRwnFN/JrF/EMeBRbzwmhG5ueiVA6
XaL1xKzFEercxAKecU2u66p8RPbmW45pFRKNm7NlYXRwjx29HT1ZIqX8RrLEQj+aosw3BQO4JmHa
4u++D05f97vR2FD+VGBmC8vZSPa1l0gK1s+ny7LdIgK0rGUvd8sR2POS8mgE5WtxHwxf/67+FTzR
8s272wYNTF4HLAEbtX7zz31rHyVQKahIspBdaKxwKc0NUlABy+GLo3JmqS5+rP1y7NbC6S3AoRx7
BZ44L/11WPAiUbRwFfSlUP78rmQSgr2+1XP5ZKeVjEBzqtmcn7EXdXFMExQfdwE5cARc63ltNn+b
AJOfC4DhHtWx5qxhYXmufYwH73dPp0Jkb+vNPFkXK2W6AJV7NnHpY5+2mq0bbS/NubHQ2pnVEj8N
QmwRWD0CZj6HQqyZ/Cv4eALjgbUsBC9iq/mM7X8c0Yw/4rNH+NgaH949+JwhUuK/8zBlMjFRneD8
P/UcPrGUFuDOZ+SEDVZH6bpwF64yFgMIl4m33EiuZTo8MrwiZdTEZFGdpafJehr6hZuwoTlBJrRp
I31edioBFaMNtZ1tvBfbmY4/wh0POLdFMEciKNxn9+VMIGeZqsSNi4ZYSjplXX6M+2f7C44Z9qo/
5Zpg+CJzv9xekHzkpBfHcuR6KERyatx5KNXrGajKu2VnhaKG8t/H+wny5NyIk9mkn9DTGBOM2QV2
mOx6uNLoTUQphmxLtcZtLxa2yF5FR28PMtF36/U1Mn+F0gqaqNS9nVD+Q/XtHGuXuFVKavLqfTYR
plfkH06DcJd5xTnbgzcnnm8Yb9MB3zOu0ZzSMPp16Dt0GLtthyIjrxpq2yByqsuKqjk68HlRO8gX
xW4KAUyBQZX2riQEB9R1Q+OsWRoYGDhvoW2oAmabe3B8gEgV2MGJrLDL68HpjnE4ZjKYUKbgMcSx
RmnOJWjwwCh/0ykzLxkLsPz8sNdw7Ts9EZve1+oP0w+K+P56ywi/XhzTHBmfvusoN+alC6r871nE
16esa72kuEbE61Nb5O92MPUd7W8u6D4rVDgArb4GfwgBKARRiAPCF5Fr4yaHZoT7i8sTk+31mGKe
KExVwq5wr6Qc9GcwEDNVvXiA5snkAQGmSQ+dyRa6lXRiM0U41Kel0VdIYYz4IutMwauIPWymPQoO
CHCtwubs38duSAC4eVDjjuhrK1ATNyJTuXLdOCljXYbw9MwCwY7A2qoy0quYg+wLuE0juaOScFWU
J4YshPRGmwhnNvt1YvW2U0CaqRAH/BAzMlk3FZISk1GdwJ6y6GOvkOs26LFrBLtSQNHAvWQt1QAn
enK7oA/+ktCNjY9c2MC4tfmvV4jpdSub62NzbamxVPEVC7fCccD7JZ1CbymrAcl1l34yKkOSxq/Z
soBn3lRNBLriL6vFHNjo/YXcvBkCmsJeJKgjL5+/KqcSqp8AvUI1C3ztbjYTyPuqrnsyB9SL78eJ
JYMYbDKtDj0gThxw+IWUaqvYI2e0GWy0IU85svxG1r4f5IctqS+pgdh9JB7YythCTEKtws3to7ib
42YKGD1Vx3g/iUmceKipLA/fbggf9T+TPE5+mmlf4k1hPI1ERhaadADPZOEhxyvwiBWZ+RBaw5yy
MAKZ9KTqbVpt6gHGw2MdxvtGrGjdmPTU8CsEHwgWqRWpWTf/CquE/elgzII940J9ArWLIk0mc/2Z
ISzI2WyRqoyFqDWiKxar7ivDqymoksNYkRNCVWEflJfqXLMs242db7hbQkwWjk7kXLdgXq+AVf02
izpmdiSOQxwIvgOuoPMb8tGSdM2A8Ox5le1ioVuu9RShgb47i9oCUIPsfFRufDxjeNDUC2lZkgCU
ZoZqdFd5NHuyEj5mM/SHJWwsPDQiP83e9w0lKRuId8Yx7cuxZJUjNQGRi98WXELCT2h9fXb/Wqss
vxV+KHb2JNO0Y3jKe9h3STYP2+CjfY8+CvuUkdNFU/CyBcIcoQJprCYtAk6zkJ1Ed6CHhSa1Ccl8
5u1lrPHu2UlrMlsGZKhyt29GUQXJ2GykvfdXMRR8wTXCKK0JiQ6UUwzFLRwivLcWxE+kRpkdcanr
DrM+05aKcmjnNIfCPyhF4Nfj/yUkom+fSnb1vDatK3uj2VbLpkQiSzM2Ty/163Al6ZeZu14afXEK
qmzGQTXUHk7rG7tuJEysFjPlsaXtkejxtrvOYgeAc2+PfNgmEQZSmVv7YS9rCEZuncNCdIhXbhsR
bYbDNWkGKUR3+4htMuB/oi0yp2SRE1wJwfKvxrrl5ahFkMVUAHCyyXldav8l1h4C7Cw1OtiDAvJz
mJE+KVScX95nzxQl0udITomPo8fs6IcblAaCuY0NbihdRFaKiHVoqu7znmKmMr30lfJKtLR/8+4U
NNNur+A7f/fUgwsOHrlySunAIrEoBi5E3uCRLF6v6ReNR0nf/QDXSdfPFv4ZnARylZ5n28pMpRz0
V2XvMN7fkXyR9oKhm5weZ/EIuPk2QeLztNDqvNbn999BEM8RIrVFsibyTHHTNoeZM7+otFFCcOLz
KoU1FMZJogFYObfDQtRdHN0ggM6fKvQIppZqPHLrDhnHS3H8h6rR/UB1xjgP4Gta9mbWNImoEij2
+CBiQS31nfePIwPZe+kC2Z5Rar8RY0vR9MoGXWKYzf50toKFi9TvQh9pDIEPYHkAlyDXTHUhqXko
j537kloP3/2W+UapTrEFxyqIhcURMqlTzNz6cd0291zo+pXad6bJNrsr+ncA8kFXumqGtttqR3b2
8TVqX/Zmi+d2h2tqXKxd0DlPfBo3cHwA16wCCzsPcmjMTsCjtLwemPj1PpWG6IclS1aySgGW8VYJ
FWcaXnbCoJZZa7khWpHrc591BHohHQfY1My9/d3OG6CM2RWBI32EJ8TGwRonvM+GKycilH8Pf1BT
ju3JkwMItAVcUX8B11vgaOc80ZPwS60U0ljhTFznAMZiLpPGWJeWrQ6yyjDZN7vT9teoCiQ8YYpq
BCRKw2bzuPsqYRVSRdfQdVnUEUrnACk3MbG0VPCGN1MSl9JNNyutswI4lIIJ5e2cY7jzQkakfATC
FluLOFJ5Ek/OYv1S7BwFkjpt3viV+OB4EbbS/m26hL+y4uzGzxkn4wnOc67CGifY7Y3uqb/tHYqR
+hB8aGcUGtCYyVe9u6vNc0HCnaq6hhnD1IZg1Jm5NjYyn+IxV9SRT3AxIn2+NsVux8Yu+c5gsAai
5v/06nybRq6NL8JkOotr2gt3V4dKa5SfFkXAOZtrSrvyoNuW34P1GyvooQGZ0LqjLvV+4ntsmwhd
2RFD9hTP7bsjF866a6wSABDBlbEfDW0FyQSAFscTFb0BeMclOaJDfoUIziB23L1LgXPjX6aJ6Hlm
ldThVoM2RDXGFFuLdWiEH552EAobtVhrBObhx80yQ+YofOyZ4zpekoHLoOcAaJ6wBEHbQGjrCIzT
4hsOsCzOZERRbygFwB+nFk/UnxR+1FvJNQXE9XauUNSWJYO55z6R4g+nThOsVMbcwG+wAozaG1v7
+b9VamVzXQONrI8RMzuZVa82nbgE7MHuZxe/jhbyyh7R7TMAyO1Ugh7HAvfyfHRj6+pj6c+hYAeV
FrY59tAqwR0AhxK4CHXcMVcyG6kS51p+hGP+YdlqP4iy/LBMK4MsUsrFo00x2b/okZ7vEJ7Q8fih
zmcgofkl9m3KLA1PQlQK4Da8H/MoC5nMXKJf8nrhSLVzT8U0USJmTaLzR++9zZxi9/tnXJSVejYn
hrusCtXYROJk3O7RbG/9gPw52x1AyJdypeRYThO/Oim3a98W11A/kG/hHGDEfouLK8PAo569O28C
cEL5Mcrf/QxhmfipNwQ25TokW4K2+eNjJiXNWRRcgd176TlnOhOmzCAGlrrII3NKSxZ92tNLgg8y
JBW/nFkukWDyey/Wyydw5mL/uTkZ6gYPU/vNs4OUMlKyUH9b5IRHmsaYHp6u54ujtCecoxjAhe7q
NCYLRMG5CCi4GIiC31qOuyACHQ1KxJAQcZ+9FSzuz5uoCFVMJKbs1hyYq5eiK3/Qt20G8w5usQPI
1VFpzTFcAXLdUvkEd8cv2wS0qsMgoWVQdII3m7THcyYpkrXNWRygYmqBhEBbr3WZePDBATyDwv3D
C7QErA5NjkGEeGjcH8/Ql4496jJtgzbXbVMAvk5s+hObTzWxBUGjwLIRm//vKOAHWlP/dPTs8WHE
tuYbKvtZ4OtvvWCkxnh/RhIOpf05Rku5J151PWVG6ej7jGkN7doyRhqH6ZoxX7tATkQXocdQsaqP
aQO2FRXJ0zHtWW17Q3owjZVuI24EPOPFThlVsIujpteXxzY/d4IC56CZ9YP+RX+EIgr/VZLdtsxb
6M3hAuP7nrp8WjYt0rKwCG1m5ougH5sI24QaSoV2vwPWnXyUIrfGrOH0iiZm/kCJxiekwZULLhya
ybUxTCjCe1YkX6BQUfkPDKu7aE6wnNl4vkOU7S6BN0YRXOUXBUtHmCymqGA+bUt75XcOn+52/n6c
ToPLc0GKbf9n8fDx7p0twQYGyRsQ0vsG5MAf5Tzynm1VkjWN8ZfqFBnoDujsFgi/DqAtbOrXj/gb
QWKNOUF2Pqp1vjeiQG/ENsQQF05rV3DAi3ZxxFZwia1AjnnwzNBlIkz0bbdjCj+wCprM8xEvWolB
OW7b7oYWmAK3C3qY3Rt/fovMP17eeTcBmpEEi0L2cRM2tqEXnCJWyX8sg0zANGUZjsvhSPVFcM9n
y/o0q5wMrmH+fdrAeeEEXzS//TyTNQTFHs9CLMfYx4iENir0b40tNp+Y3YrcO+TALJiJiWQLCoqU
RixiaHCeSkLMx88EuZk/puhVcLhaY9epqRskulr4JV+vBxcD+iuYHrqlzmRskAinoFQr91pajvPw
xNyydrTFlQhlZKEocOwOsLoXgKzZImAytHRJrf0dcvLMzsNLTETlIvEE8VS22vwsbGDAxb+yKnOn
67qiNmz/de66OFHwoutYbbkXytBuGOzYzI1Ku5gRxZjnJYvm1Vw8dDDlVq3yQYEJp885nAmvpeya
2G/yLdh7flp5WbE9rJh4bWqDYg2OJ6gRlIfYwgK7e8BYohlWlhCB9nWBMzO0uF57h+z906GpqYLF
tajxvIuiLc36PpMdbTCOSVaUKAd4R/bUXjSutXWwNoUf5o9y38m+phTLSeD5aUtvgRv1YXaHOar9
vduJeMV7/OsqDBXHTKzTCk1EHl0qSSdaf7mG9kRPnB92EXlwUKWWDwAxS4B6/Q82XbCx38cQN3GI
3gMTwdRV8IRb65ohhG/yURQ5AxaNk3HZI+80/zuC0gdId/q1NV+TNNJz79E9uQRrn3y9N9hrnUk8
S5iBUJI7RWcgooMSIa5buG5I0MRXVafjdB8kNukSCiu0u2bwkE4MDcDbLEdYssWc+CAzVjafKEu3
rham2O47CxIDzpow3aKG3WkU1aaiMPKgpE/ZjrS4cj/4RMuyMp1WvGc6dUEjEUnww/tTF3ut5BYX
xkIufjk8po4J3r6rurTc27YjYIFHbLZjtwbofPBca3fXPxCOaQfjaJpsfCs1M2qtrCZqC8XQzqtL
b0nyZ2QZM0aTOdXfjeS/rylOxgFG4Vpyc8CW34+jWeMNY35vJyi0H3nz+fCtFH+OX/nzOrMdjhtA
D3ZUIibtmPPTvc6BFfiDbYY0wW8OIM9LK38io3asqiRGG697XEvgX8nFSM4mGJk8JmXHhsSbE4su
QpQxx/LW0063etHPpIKs2EBh122uxtyklYHb/TVOk5L4tloRhgMCgNjw44RdpK8PbsdHBEbuNyLE
ANT1teJuL/mhRPA18f8x8qzROZVEfIIYnBfqx5e36GG30S32s24XhwPCjDKsX384bXDhZ2LCzbq+
pUB/GOtVAAzGkPanv4+FmR7y9tYBMfczbRlvyNcyN7upK1WVsTCI+Wb93gYm9AJYj5dwtJxvLQV+
jUaJhpfge8NQpjlUhmOecG1zFqyBecd4nbVzUhpKmFvMyYv/5BR7txHXT1ljyc/nueg8H8EL2tUH
qDOo0aMXdoyzoBkkkHcWYGFVxBuYgJrjYeYT/MQ1crOnA6ummbEcCM5gN9h1CRCHMfLU2X/BqUwk
QG0LXLNDC0sFLq0MSIyghjNtoLfdXUuquMVnrBuqZ+ScYCl84Blhd2yL8NPdsemOk2WifOSJMIMf
XqSRqsEZXyZ//CTdmpilMJj4lOSAGttJkyuGnKcpz8dOvYQmkuWxmUWlO0oQAmVoq3jdxGOoQoMY
y9I44jH3NahcCK3Qoen+SRSVM6BDCCrYMwq7Boqn11E9qMS8iDDrIiQhiBehmU3OX9nMI7MC7Ld/
N31XyjPBjCmdtdRxHgMkbSBlNN53xGzonxNUTp75c8CUzAkYrR/kZGfdWkavUVa19g4dpcDxQWR/
uuE4VT8R+7o9A5CWOGOJpgeVgqWXz/m54KLhaOWG6JjNZXwnUfQc5+Ux5Ip4tfIS4PnKM8anIEwc
Cd0lR0jgGBIj2kDo1epmVn71hchshCVJmSRwv18BbtJiWmTBEySCQqelQk2qyiFk1RvB3hp1TD4x
Z378wXmrnYa40uUGqvTjySeodfdWMun89uIh8uNaDmlS+mcyGdNq6KOVkFtS/LXWFRVgqIkbnuyL
JlKkuIeiFjWbEIdtdwByE6dHN6FAFUg0GQeLHqJ7FWH6kaVRpYO0NDAtX7byVWHYvVVVein3VB2g
my2MPpW0eZT0oMOYUy5ubzQbIJHk6nc+rmz1wNrBkytmbOtW77ZvUi+2595229KZEHltEEfBjOEY
1nbXavZ1jxlEGnPjdQeUya4PPFOZfwts16U36me9nVo4Feo+6mpZpdmFC1EAP/ELhMEU2lqbhoYV
aKBdB8NMsCagNA6H071aSZpGJtWiBqPAB3NokECeHPSVGjuBU3JWpDxMQEd4c2IKQqi1jCO/ZMNM
MGEcQp4yUojI0UQyH953SfhaXDssdrLjI78mXKXUxGAvZ3gL9b4DsBQbPddBKRwRZEOGlf1w7jSB
IzKJIW8kb18zLzK5ITWn2yI1RyVaeDvuE0oN3+I6VWIC+cXEwFKccLtau0eDQM3KKO1bMHyqUz2q
KhLDASL7K9lWS2sFxur+03nfldLD4QoSx+2Q5fQ0zYczBTX1kZEQ++9a5wYnSXJhB7h6FGqSXn7t
wvRoQtrI96/Thj3hd1npuA==
`protect end_protected
